module ProcessamentoDigito(
	input  [7:0] numero[10:0][10:0],
	input flag,
	output [3:0] digito
);
	
	wire [15:0] v_diferenca[9:0];
	wire [7:0] diff_pixel[9:0][10:0][10:0];
	
	SomaPixels somaPixels0(diff_pixel[0],flag,v_diferenca[0]);
	SomaPixels somaPixels1(diff_pixel[1],flag,v_diferenca[1]);
	SomaPixels somaPixels2(diff_pixel[2],flag,v_diferenca[2]);
	SomaPixels somaPixels3(diff_pixel[3],flag,v_diferenca[3]);
	SomaPixels somaPixels4(diff_pixel[4],flag,v_diferenca[4]);
	SomaPixels somaPixels5(diff_pixel[5],flag,v_diferenca[5]);
	SomaPixels somaPixels6(diff_pixel[6],flag,v_diferenca[6]);
	SomaPixels somaPixels7(diff_pixel[7],flag,v_diferenca[7]);
	SomaPixels somaPixels8(diff_pixel[8],flag,v_diferenca[8]);
	SomaPixels somaPixels9(diff_pixel[9],flag,v_diferenca[9]);
	
	MenorDistancia menorDistancia(v_diferenca, flag, digito);
	
	always@(posedge flag)
	begin
	
		//diff_pixel[00][00][00] <= numero[00][00] > 26 ? numero[00][00] - 26 : 26 - numero[00][00];
		//diff_pixel[00][00][01] <= numero[00][01] > 27 ? numero[00][01] - 27 : 27 - numero[00][01];
		//diff_pixel[00][00][02] <= numero[00][02] > 37 ? numero[00][02] - 37 : 37 - numero[00][02];
		//diff_pixel[00][00][03] <= numero[00][03] > 67 ? numero[00][03] - 67 : 67 - numero[00][03];
		//diff_pixel[00][00][04] <= numero[00][04] > 86 ? numero[00][04] - 86 : 86 - numero[00][04];
		//diff_pixel[00][00][05] <= numero[00][05] > 97 ? numero[00][05] - 97 : 97 - numero[00][05];
		//diff_pixel[00][00][06] <= numero[00][06] > 86 ? numero[00][06] - 86 : 86 - numero[00][06];
		//diff_pixel[00][00][07] <= numero[00][07] > 64 ? numero[00][07] - 64 : 64 - numero[00][07];
		//diff_pixel[00][00][08] <= numero[00][08] > 27 ? numero[00][08] - 27 : 27 - numero[00][08];
		//diff_pixel[00][00][09] <= numero[00][09] > 5 ? numero[00][09] - 5 : 5 - numero[00][09];
		//diff_pixel[00][00][10] <= numero[00][10] > 0 ? numero[00][10] - 0 : 0 - numero[00][10];
		//diff_pixel[00][01][00] <= numero[01][00] > 17 ? numero[01][00] - 17 : 17 - numero[01][00];
		//diff_pixel[00][01][01] <= numero[01][01] > 28 ? numero[01][01] - 28 : 28 - numero[01][01];
		//diff_pixel[00][01][02] <= numero[01][02] > 57 ? numero[01][02] - 57 : 57 - numero[01][02];
		//diff_pixel[00][01][03] <= numero[01][03] > 93 ? numero[01][03] - 93 : 93 - numero[01][03];
		//diff_pixel[00][01][04] <= numero[01][04] > 123 ? numero[01][04] - 123 : 123 - numero[01][04];
		//diff_pixel[00][01][05] <= numero[01][05] > 138 ? numero[01][05] - 138 : 138 - numero[01][05];
		//diff_pixel[00][01][06] <= numero[01][06] > 135 ? numero[01][06] - 135 : 135 - numero[01][06];
		//diff_pixel[00][01][07] <= numero[01][07] > 116 ? numero[01][07] - 116 : 116 - numero[01][07];
		//diff_pixel[00][01][08] <= numero[01][08] > 74 ? numero[01][08] - 74 : 74 - numero[01][08];
		//diff_pixel[00][01][09] <= numero[01][09] > 36 ? numero[01][09] - 36 : 36 - numero[01][09];
		//diff_pixel[00][01][10] <= numero[01][10] > 7 ? numero[01][10] - 7 : 7 - numero[01][10];
		diff_pixel[00][02][00] <= numero[02][00] > 23 ? numero[02][00] - 23 : 23 - numero[02][00];
		diff_pixel[00][02][01] <= numero[02][01] > 51 ? numero[02][01] - 51 : 51 - numero[02][01];
		diff_pixel[00][02][02] <= numero[02][02] > 75 ? numero[02][02] - 75 : 75 - numero[02][02];
		diff_pixel[00][02][03] <= numero[02][03] > 63 ? numero[02][03] - 63 : 63 - numero[02][03];
		diff_pixel[00][02][04] <= numero[02][04] > 58 ? numero[02][04] - 58 : 58 - numero[02][04];
		diff_pixel[00][02][05] <= numero[02][05] > 63 ? numero[02][05] - 63 : 63 - numero[02][05];
		diff_pixel[00][02][06] <= numero[02][06] > 91 ? numero[02][06] - 91 : 91 - numero[02][06];
		diff_pixel[00][02][07] <= numero[02][07] > 123 ? numero[02][07] - 123 : 123 - numero[02][07];
		diff_pixel[00][02][08] <= numero[02][08] > 125 ? numero[02][08] - 125 : 125 - numero[02][08];
		diff_pixel[00][02][09] <= numero[02][09] > 95 ? numero[02][09] - 95 : 95 - numero[02][09];
		diff_pixel[00][02][10] <= numero[02][10] > 45 ? numero[02][10] - 45 : 45 - numero[02][10];
		diff_pixel[00][03][00] <= numero[03][00] > 77 ? numero[03][00] - 77 : 77 - numero[03][00];
		diff_pixel[00][03][01] <= numero[03][01] > 101 ? numero[03][01] - 101 : 101 - numero[03][01];
		diff_pixel[00][03][02] <= numero[03][02] > 103 ? numero[03][02] - 103 : 103 - numero[03][02];
		diff_pixel[00][03][03] <= numero[03][03] > 69 ? numero[03][03] - 69 : 69 - numero[03][03];
		diff_pixel[00][03][04] <= numero[03][04] > 34 ? numero[03][04] - 34 : 34 - numero[03][04];
		diff_pixel[00][03][05] <= numero[03][05] > 23 ? numero[03][05] - 23 : 23 - numero[03][05];
		diff_pixel[00][03][06] <= numero[03][06] > 44 ? numero[03][06] - 44 : 44 - numero[03][06];
		diff_pixel[00][03][07] <= numero[03][07] > 81 ? numero[03][07] - 81 : 81 - numero[03][07];
		diff_pixel[00][03][08] <= numero[03][08] > 113 ? numero[03][08] - 113 : 113 - numero[03][08];
		diff_pixel[00][03][09] <= numero[03][09] > 111 ? numero[03][09] - 111 : 111 - numero[03][09];
		diff_pixel[00][03][10] <= numero[03][10] > 92 ? numero[03][10] - 92 : 92 - numero[03][10];
		diff_pixel[00][04][00] <= numero[04][00] > 105 ? numero[04][00] - 105 : 105 - numero[04][00];
		diff_pixel[00][04][01] <= numero[04][01] > 129 ? numero[04][01] - 129 : 129 - numero[04][01];
		diff_pixel[00][04][02] <= numero[04][02] > 123 ? numero[04][02] - 123 : 123 - numero[04][02];
		diff_pixel[00][04][03] <= numero[04][03] > 81 ? numero[04][03] - 81 : 81 - numero[04][03];
		diff_pixel[00][04][04] <= numero[04][04] > 36 ? numero[04][04] - 36 : 36 - numero[04][04];
		diff_pixel[00][04][05] <= numero[04][05] > 12 ? numero[04][05] - 12 : 12 - numero[04][05];
		diff_pixel[00][04][06] <= numero[04][06] > 26 ? numero[04][06] - 26 : 26 - numero[04][06];
		diff_pixel[00][04][07] <= numero[04][07] > 66 ? numero[04][07] - 66 : 66 - numero[04][07];
		diff_pixel[00][04][08] <= numero[04][08] > 117 ? numero[04][08] - 117 : 117 - numero[04][08];
		diff_pixel[00][04][09] <= numero[04][09] > 133 ? numero[04][09] - 133 : 133 - numero[04][09];
		diff_pixel[00][04][10] <= numero[04][10] > 129 ? numero[04][10] - 129 : 129 - numero[04][10];
		diff_pixel[00][05][00] <= numero[05][00] > 105 ? numero[05][00] - 105 : 105 - numero[05][00];
		diff_pixel[00][05][01] <= numero[05][01] > 129 ? numero[05][01] - 129 : 129 - numero[05][01];
		diff_pixel[00][05][02] <= numero[05][02] > 122 ? numero[05][02] - 122 : 122 - numero[05][02];
		diff_pixel[00][05][03] <= numero[05][03] > 80 ? numero[05][03] - 80 : 80 - numero[05][03];
		diff_pixel[00][05][04] <= numero[05][04] > 30 ? numero[05][04] - 30 : 30 - numero[05][04];
		diff_pixel[00][05][05] <= numero[05][05] > 8 ? numero[05][05] - 8 : 8 - numero[05][05];
		diff_pixel[00][05][06] <= numero[05][06] > 22 ? numero[05][06] - 22 : 22 - numero[05][06];
		diff_pixel[00][05][07] <= numero[05][07] > 62 ? numero[05][07] - 62 : 62 - numero[05][07];
		diff_pixel[00][05][08] <= numero[05][08] > 111 ? numero[05][08] - 111 : 111 - numero[05][08];
		diff_pixel[00][05][09] <= numero[05][09] > 126 ? numero[05][09] - 126 : 126 - numero[05][09];
		diff_pixel[00][05][10] <= numero[05][10] > 125 ? numero[05][10] - 125 : 125 - numero[05][10];
		diff_pixel[00][06][00] <= numero[06][00] > 112 ? numero[06][00] - 112 : 112 - numero[06][00];
		diff_pixel[00][06][01] <= numero[06][01] > 123 ? numero[06][01] - 123 : 123 - numero[06][01];
		diff_pixel[00][06][02] <= numero[06][02] > 116 ? numero[06][02] - 116 : 116 - numero[06][02];
		diff_pixel[00][06][03] <= numero[06][03] > 76 ? numero[06][03] - 76 : 76 - numero[06][03];
		diff_pixel[00][06][04] <= numero[06][04] > 28 ? numero[06][04] - 28 : 28 - numero[06][04];
		diff_pixel[00][06][05] <= numero[06][05] > 4 ? numero[06][05] - 4 : 4 - numero[06][05];
		diff_pixel[00][06][06] <= numero[06][06] > 19 ? numero[06][06] - 19 : 19 - numero[06][06];
		diff_pixel[00][06][07] <= numero[06][07] > 59 ? numero[06][07] - 59 : 59 - numero[06][07];
		diff_pixel[00][06][08] <= numero[06][08] > 110 ? numero[06][08] - 110 : 110 - numero[06][08];
		diff_pixel[00][06][09] <= numero[06][09] > 126 ? numero[06][09] - 126 : 126 - numero[06][09];
		diff_pixel[00][06][10] <= numero[06][10] > 125 ? numero[06][10] - 125 : 125 - numero[06][10];
		diff_pixel[00][07][00] <= numero[07][00] > 97 ? numero[07][00] - 97 : 97 - numero[07][00];
		diff_pixel[00][07][01] <= numero[07][01] > 108 ? numero[07][01] - 108 : 108 - numero[07][01];
		diff_pixel[00][07][02] <= numero[07][02] > 116 ? numero[07][02] - 116 : 116 - numero[07][02];
		diff_pixel[00][07][03] <= numero[07][03] > 93 ? numero[07][03] - 93 : 93 - numero[07][03];
		diff_pixel[00][07][04] <= numero[07][04] > 54 ? numero[07][04] - 54 : 54 - numero[07][04];
		diff_pixel[00][07][05] <= numero[07][05] > 23 ? numero[07][05] - 23 : 23 - numero[07][05];
		diff_pixel[00][07][06] <= numero[07][06] > 27 ? numero[07][06] - 27 : 27 - numero[07][06];
		diff_pixel[00][07][07] <= numero[07][07] > 56 ? numero[07][07] - 56 : 56 - numero[07][07];
		diff_pixel[00][07][08] <= numero[07][08] > 97 ? numero[07][08] - 97 : 97 - numero[07][08];
		diff_pixel[00][07][09] <= numero[07][09] > 110 ? numero[07][09] - 110 : 110 - numero[07][09];
		diff_pixel[00][07][10] <= numero[07][10] > 97 ? numero[07][10] - 97 : 97 - numero[07][10];
		//diff_pixel[00][08][00] <= numero[08][00] > 42 ? numero[08][00] - 42 : 42 - numero[08][00];
		//diff_pixel[00][08][01] <= numero[08][01] > 71 ? numero[08][01] - 71 : 71 - numero[08][01];
		//diff_pixel[00][08][02] <= numero[08][02] > 109 ? numero[08][02] - 109 : 109 - numero[08][02];
		//diff_pixel[00][08][03] <= numero[08][03] > 121 ? numero[08][03] - 121 : 121 - numero[08][03];
		//diff_pixel[00][08][04] <= numero[08][04] > 94 ? numero[08][04] - 94 : 94 - numero[08][04];
		//diff_pixel[00][08][05] <= numero[08][05] > 49 ? numero[08][05] - 49 : 49 - numero[08][05];
		//diff_pixel[00][08][06] <= numero[08][06] > 39 ? numero[08][06] - 39 : 39 - numero[08][06];
		//diff_pixel[00][08][07] <= numero[08][07] > 40 ? numero[08][07] - 40 : 40 - numero[08][07];
		//diff_pixel[00][08][08] <= numero[08][08] > 67 ? numero[08][08] - 67 : 67 - numero[08][08];
		//diff_pixel[00][08][09] <= numero[08][09] > 65 ? numero[08][09] - 65 : 65 - numero[08][09];
		//diff_pixel[00][08][10] <= numero[08][10] > 41 ? numero[08][10] - 41 : 41 - numero[08][10];
		//diff_pixel[00][09][00] <= numero[09][00] > 5 ? numero[09][00] - 5 : 5 - numero[09][00];
		//diff_pixel[00][09][01] <= numero[09][01] > 30 ? numero[09][01] - 30 : 30 - numero[09][01];
		//diff_pixel[00][09][02] <= numero[09][02] > 70 ? numero[09][02] - 70 : 70 - numero[09][02];
		//diff_pixel[00][09][03] <= numero[09][03] > 108 ? numero[09][03] - 108 : 108 - numero[09][03];
		//diff_pixel[00][09][04] <= numero[09][04] > 131 ? numero[09][04] - 131 : 131 - numero[09][04];
		//diff_pixel[00][09][05] <= numero[09][05] > 131 ? numero[09][05] - 131 : 131 - numero[09][05];
		//diff_pixel[00][09][06] <= numero[09][06] > 115 ? numero[09][06] - 115 : 115 - numero[09][06];
		//diff_pixel[00][09][07] <= numero[09][07] > 90 ? numero[09][07] - 90 : 90 - numero[09][07];
		//diff_pixel[00][09][08] <= numero[09][08] > 57 ? numero[09][08] - 57 : 57 - numero[09][08];
		//diff_pixel[00][09][09] <= numero[09][09] > 30 ? numero[09][09] - 30 : 30 - numero[09][09];
		//diff_pixel[00][09][10] <= numero[09][10] > 7 ? numero[09][10] - 7 : 7 - numero[09][10];
		//diff_pixel[00][10][00] <= numero[10][00] > 0 ? numero[10][00] - 0 : 0 - numero[10][00];
		//diff_pixel[00][10][01] <= numero[10][01] > 7 ? numero[10][01] - 7 : 7 - numero[10][01];
		//diff_pixel[00][10][02] <= numero[10][02] > 28 ? numero[10][02] - 28 : 28 - numero[10][02];
		//diff_pixel[00][10][03] <= numero[10][03] > 62 ? numero[10][03] - 62 : 62 - numero[10][03];
		//diff_pixel[00][10][04] <= numero[10][04] > 90 ? numero[10][04] - 90 : 90 - numero[10][04];
		//diff_pixel[00][10][05] <= numero[10][05] > 104 ? numero[10][05] - 104 : 104 - numero[10][05];
		//diff_pixel[00][10][06] <= numero[10][06] > 99 ? numero[10][06] - 99 : 99 - numero[10][06];
		//diff_pixel[00][10][07] <= numero[10][07] > 73 ? numero[10][07] - 73 : 73 - numero[10][07];
		//diff_pixel[00][10][08] <= numero[10][08] > 39 ? numero[10][08] - 39 : 39 - numero[10][08];
		//diff_pixel[00][10][09] <= numero[10][09] > 11 ? numero[10][09] - 11 : 11 - numero[10][09];
		//diff_pixel[00][10][10] <= numero[10][10] > 0 ? numero[10][10] - 0 : 0 - numero[10][10];
		
		//diff_pixel[01][00][00] <= numero[00][00] > 0 ? numero[00][00] - 0 : 0 - numero[00][00];
		//diff_pixel[01][00][01] <= numero[00][01] > 0 ? numero[00][01] - 0 : 0 - numero[00][01];
		//diff_pixel[01][00][02] <= numero[00][02] > 0 ? numero[00][02] - 0 : 0 - numero[00][02];
		//diff_pixel[01][00][03] <= numero[00][03] > 12 ? numero[00][03] - 12 : 12 - numero[00][03];
		//diff_pixel[01][00][04] <= numero[00][04] > 36 ? numero[00][04] - 36 : 36 - numero[00][04];
		//diff_pixel[01][00][05] <= numero[00][05] > 62 ? numero[00][05] - 62 : 62 - numero[00][05];
		//diff_pixel[01][00][06] <= numero[00][06] > 69 ? numero[00][06] - 69 : 69 - numero[00][06];
		//diff_pixel[01][00][07] <= numero[00][07] > 60 ? numero[00][07] - 60 : 60 - numero[00][07];
		//diff_pixel[01][00][08] <= numero[00][08] > 35 ? numero[00][08] - 35 : 35 - numero[00][08];
		//diff_pixel[01][00][09] <= numero[00][09] > 9 ? numero[00][09] - 9 : 9 - numero[00][09];
		//diff_pixel[01][00][10] <= numero[00][10] > 0 ? numero[00][10] - 0 : 0 - numero[00][10];
		//diff_pixel[01][01][00] <= numero[01][00] > 0 ? numero[01][00] - 0 : 0 - numero[01][00];
		//diff_pixel[01][01][01] <= numero[01][01] > 0 ? numero[01][01] - 0 : 0 - numero[01][01];
		//diff_pixel[01][01][02] <= numero[01][02] > 13 ? numero[01][02] - 13 : 13 - numero[01][02];
		//diff_pixel[01][01][03] <= numero[01][03] > 46 ? numero[01][03] - 46 : 46 - numero[01][03];
		//diff_pixel[01][01][04] <= numero[01][04] > 88 ? numero[01][04] - 88 : 88 - numero[01][04];
		//diff_pixel[01][01][05] <= numero[01][05] > 128 ? numero[01][05] - 128 : 128 - numero[01][05];
		//diff_pixel[01][01][06] <= numero[01][06] > 136 ? numero[01][06] - 136 : 136 - numero[01][06];
		//diff_pixel[01][01][07] <= numero[01][07] > 113 ? numero[01][07] - 113 : 113 - numero[01][07];
		//diff_pixel[01][01][08] <= numero[01][08] > 65 ? numero[01][08] - 65 : 65 - numero[01][08];
		//diff_pixel[01][01][09] <= numero[01][09] > 22 ? numero[01][09] - 22 : 22 - numero[01][09];
		//diff_pixel[01][01][10] <= numero[01][10] > 0 ? numero[01][10] - 0 : 0 - numero[01][10];
		diff_pixel[01][02][00] <= numero[02][00] > 0 ? numero[02][00] - 0 : 0 - numero[02][00];
		diff_pixel[01][02][01] <= numero[02][01] > 11 ? numero[02][01] - 11 : 11 - numero[02][01];
		diff_pixel[01][02][02] <= numero[02][02] > 47 ? numero[02][02] - 47 : 47 - numero[02][02];
		diff_pixel[01][02][03] <= numero[02][03] > 95 ? numero[02][03] - 95 : 95 - numero[02][03];
		diff_pixel[01][02][04] <= numero[02][04] > 143 ? numero[02][04] - 143 : 143 - numero[02][04];
		diff_pixel[01][02][05] <= numero[02][05] > 167 ? numero[02][05] - 167 : 167 - numero[02][05];
		diff_pixel[01][02][06] <= numero[02][06] > 154 ? numero[02][06] - 154 : 154 - numero[02][06];
		diff_pixel[01][02][07] <= numero[02][07] > 118 ? numero[02][07] - 118 : 118 - numero[02][07];
		diff_pixel[01][02][08] <= numero[02][08] > 60 ? numero[02][08] - 60 : 60 - numero[02][08];
		diff_pixel[01][02][09] <= numero[02][09] > 19 ? numero[02][09] - 19 : 19 - numero[02][09];
		diff_pixel[01][02][10] <= numero[02][10] > 0 ? numero[02][10] - 0 : 0 - numero[02][10];
		diff_pixel[01][03][00] <= numero[03][00] > 1 ? numero[03][00] - 1 : 1 - numero[03][00];
		diff_pixel[01][03][01] <= numero[03][01] > 0 ? numero[03][01] - 0 : 0 - numero[03][01];
		diff_pixel[01][03][02] <= numero[03][02] > 18 ? numero[03][02] - 18 : 18 - numero[03][02];
		diff_pixel[01][03][03] <= numero[03][03] > 56 ? numero[03][03] - 56 : 56 - numero[03][03];
		diff_pixel[01][03][04] <= numero[03][04] > 99 ? numero[03][04] - 99 : 99 - numero[03][04];
		diff_pixel[01][03][05] <= numero[03][05] > 137 ? numero[03][05] - 137 : 137 - numero[03][05];
		diff_pixel[01][03][06] <= numero[03][06] > 139 ? numero[03][06] - 139 : 139 - numero[03][06];
		diff_pixel[01][03][07] <= numero[03][07] > 115 ? numero[03][07] - 115 : 115 - numero[03][07];
		diff_pixel[01][03][08] <= numero[03][08] > 62 ? numero[03][08] - 62 : 62 - numero[03][08];
		diff_pixel[01][03][09] <= numero[03][09] > 19 ? numero[03][09] - 19 : 19 - numero[03][09];
		diff_pixel[01][03][10] <= numero[03][10] > 3 ? numero[03][10] - 3 : 3 - numero[03][10];
		diff_pixel[01][04][00] <= numero[04][00] > 1 ? numero[04][00] - 1 : 1 - numero[04][00];
		diff_pixel[01][04][01] <= numero[04][01] > 0 ? numero[04][01] - 0 : 0 - numero[04][01];
		diff_pixel[01][04][02] <= numero[04][02] > 0 ? numero[04][02] - 0 : 0 - numero[04][02];
		diff_pixel[01][04][03] <= numero[04][03] > 26 ? numero[04][03] - 26 : 26 - numero[04][03];
		diff_pixel[01][04][04] <= numero[04][04] > 71 ? numero[04][04] - 71 : 71 - numero[04][04];
		diff_pixel[01][04][05] <= numero[04][05] > 117 ? numero[04][05] - 117 : 117 - numero[04][05];
		diff_pixel[01][04][06] <= numero[04][06] > 129 ? numero[04][06] - 129 : 129 - numero[04][06];
		diff_pixel[01][04][07] <= numero[04][07] > 112 ? numero[04][07] - 112 : 112 - numero[04][07];
		diff_pixel[01][04][08] <= numero[04][08] > 64 ? numero[04][08] - 64 : 64 - numero[04][08];
		diff_pixel[01][04][09] <= numero[04][09] > 17 ? numero[04][09] - 17 : 17 - numero[04][09];
		diff_pixel[01][04][10] <= numero[04][10] > 2 ? numero[04][10] - 2 : 2 - numero[04][10];
		diff_pixel[01][05][00] <= numero[05][00] > 5 ? numero[05][00] - 5 : 5 - numero[05][00];
		diff_pixel[01][05][01] <= numero[05][01] > 0 ? numero[05][01] - 0 : 0 - numero[05][01];
		diff_pixel[01][05][02] <= numero[05][02] > 0 ? numero[05][02] - 0 : 0 - numero[05][02];
		diff_pixel[01][05][03] <= numero[05][03] > 28 ? numero[05][03] - 28 : 28 - numero[05][03];
		diff_pixel[01][05][04] <= numero[05][04] > 71 ? numero[05][04] - 71 : 71 - numero[05][04];
		diff_pixel[01][05][05] <= numero[05][05] > 117 ? numero[05][05] - 117 : 117 - numero[05][05];
		diff_pixel[01][05][06] <= numero[05][06] > 129 ? numero[05][06] - 129 : 129 - numero[05][06];
		diff_pixel[01][05][07] <= numero[05][07] > 112 ? numero[05][07] - 112 : 112 - numero[05][07];
		diff_pixel[01][05][08] <= numero[05][08] > 63 ? numero[05][08] - 63 : 63 - numero[05][08];
		diff_pixel[01][05][09] <= numero[05][09] > 17 ? numero[05][09] - 17 : 17 - numero[05][09];
		diff_pixel[01][05][10] <= numero[05][10] > 4 ? numero[05][10] - 4 : 4 - numero[05][10];
		diff_pixel[01][06][00] <= numero[06][00] > 6 ? numero[06][00] - 6 : 6 - numero[06][00];
		diff_pixel[01][06][01] <= numero[06][01] > 0 ? numero[06][01] - 0 : 0 - numero[06][01];
		diff_pixel[01][06][02] <= numero[06][02] > 0 ? numero[06][02] - 0 : 0 - numero[06][02];
		diff_pixel[01][06][03] <= numero[06][03] > 29 ? numero[06][03] - 29 : 29 - numero[06][03];
		diff_pixel[01][06][04] <= numero[06][04] > 70 ? numero[06][04] - 70 : 70 - numero[06][04];
		diff_pixel[01][06][05] <= numero[06][05] > 116 ? numero[06][05] - 116 : 116 - numero[06][05];
		diff_pixel[01][06][06] <= numero[06][06] > 128 ? numero[06][06] - 128 : 128 - numero[06][06];
		diff_pixel[01][06][07] <= numero[06][07] > 111 ? numero[06][07] - 111 : 111 - numero[06][07];
		diff_pixel[01][06][08] <= numero[06][08] > 63 ? numero[06][08] - 63 : 63 - numero[06][08];
		diff_pixel[01][06][09] <= numero[06][09] > 16 ? numero[06][09] - 16 : 16 - numero[06][09];
		diff_pixel[01][06][10] <= numero[06][10] > 5 ? numero[06][10] - 5 : 5 - numero[06][10];
		diff_pixel[01][07][00] <= numero[07][00] > 2 ? numero[07][00] - 2 : 2 - numero[07][00];
		diff_pixel[01][07][01] <= numero[07][01] > 0 ? numero[07][01] - 0 : 0 - numero[07][01];
		diff_pixel[01][07][02] <= numero[07][02] > 0 ? numero[07][02] - 0 : 0 - numero[07][02];
		diff_pixel[01][07][03] <= numero[07][03] > 29 ? numero[07][03] - 29 : 29 - numero[07][03];
		diff_pixel[01][07][04] <= numero[07][04] > 71 ? numero[07][04] - 71 : 71 - numero[07][04];
		diff_pixel[01][07][05] <= numero[07][05] > 117 ? numero[07][05] - 117 : 117 - numero[07][05];
		diff_pixel[01][07][06] <= numero[07][06] > 128 ? numero[07][06] - 128 : 128 - numero[07][06];
		diff_pixel[01][07][07] <= numero[07][07] > 113 ? numero[07][07] - 113 : 113 - numero[07][07];
		diff_pixel[01][07][08] <= numero[07][08] > 61 ? numero[07][08] - 61 : 61 - numero[07][08];
		diff_pixel[01][07][09] <= numero[07][09] > 15 ? numero[07][09] - 15 : 15 - numero[07][09];
		diff_pixel[01][07][10] <= numero[07][10] > 1 ? numero[07][10] - 1 : 1 - numero[07][10];
		//diff_pixel[01][08][00] <= numero[08][00] > 0 ? numero[08][00] - 0 : 0 - numero[08][00];
		//diff_pixel[01][08][01] <= numero[08][01] > 0 ? numero[08][01] - 0 : 0 - numero[08][01];
		//diff_pixel[01][08][02] <= numero[08][02] > 2 ? numero[08][02] - 2 : 2 - numero[08][02];
		//diff_pixel[01][08][03] <= numero[08][03] > 29 ? numero[08][03] - 29 : 29 - numero[08][03];
		//diff_pixel[01][08][04] <= numero[08][04] > 68 ? numero[08][04] - 68 : 68 - numero[08][04];
		//diff_pixel[01][08][05] <= numero[08][05] > 116 ? numero[08][05] - 116 : 116 - numero[08][05];
		//diff_pixel[01][08][06] <= numero[08][06] > 131 ? numero[08][06] - 131 : 131 - numero[08][06];
		//diff_pixel[01][08][07] <= numero[08][07] > 115 ? numero[08][07] - 115 : 115 - numero[08][07];
		//diff_pixel[01][08][08] <= numero[08][08] > 69 ? numero[08][08] - 69 : 69 - numero[08][08];
		//diff_pixel[01][08][09] <= numero[08][09] > 24 ? numero[08][09] - 24 : 24 - numero[08][09];
		//diff_pixel[01][08][10] <= numero[08][10] > 1 ? numero[08][10] - 1 : 1 - numero[08][10];
		//diff_pixel[01][09][00] <= numero[09][00] > 22 ? numero[09][00] - 22 : 22 - numero[09][00];
		//diff_pixel[01][09][01] <= numero[09][01] > 54 ? numero[09][01] - 54 : 54 - numero[09][01];
		//diff_pixel[01][09][02] <= numero[09][02] > 93 ? numero[09][02] - 93 : 93 - numero[09][02];
		//diff_pixel[01][09][03] <= numero[09][03] > 125 ? numero[09][03] - 125 : 125 - numero[09][03];
		//diff_pixel[01][09][04] <= numero[09][04] > 149 ? numero[09][04] - 149 : 149 - numero[09][04];
		//diff_pixel[01][09][05] <= numero[09][05] > 165 ? numero[09][05] - 165 : 165 - numero[09][05];
		//diff_pixel[01][09][06] <= numero[09][06] > 165 ? numero[09][06] - 165 : 165 - numero[09][06];
		//diff_pixel[01][09][07] <= numero[09][07] > 159 ? numero[09][07] - 159 : 159 - numero[09][07];
		//diff_pixel[01][09][08] <= numero[09][08] > 139 ? numero[09][08] - 139 : 139 - numero[09][08];
		//diff_pixel[01][09][09] <= numero[09][09] > 109 ? numero[09][09] - 109 : 109 - numero[09][09];
		//diff_pixel[01][09][10] <= numero[09][10] > 79 ? numero[09][10] - 79 : 79 - numero[09][10];
		//diff_pixel[01][10][00] <= numero[10][00] > 15 ? numero[10][00] - 15 : 15 - numero[10][00];
		//diff_pixel[01][10][01] <= numero[10][01] > 46 ? numero[10][01] - 46 : 46 - numero[10][01];
		//diff_pixel[01][10][02] <= numero[10][02] > 82 ? numero[10][02] - 82 : 82 - numero[10][02];
		//diff_pixel[01][10][03] <= numero[10][03] > 106 ? numero[10][03] - 106 : 106 - numero[10][03];
		//diff_pixel[01][10][04] <= numero[10][04] > 118 ? numero[10][04] - 118 : 118 - numero[10][04];
		//diff_pixel[01][10][05] <= numero[10][05] > 120 ? numero[10][05] - 120 : 120 - numero[10][05];
		//diff_pixel[01][10][06] <= numero[10][06] > 122 ? numero[10][06] - 122 : 122 - numero[10][06];
		//diff_pixel[01][10][07] <= numero[10][07] > 122 ? numero[10][07] - 122 : 122 - numero[10][07];
		//diff_pixel[01][10][08] <= numero[10][08] > 122 ? numero[10][08] - 122 : 122 - numero[10][08];
		//diff_pixel[01][10][09] <= numero[10][09] > 107 ? numero[10][09] - 107 : 107 - numero[10][09];
		//diff_pixel[01][10][10] <= numero[10][10] > 82 ? numero[10][10] - 82 : 82 - numero[10][10];
		
		//diff_pixel[02][00][00] <= numero[00][00] > 30 ? numero[00][00] - 30 : 30 - numero[00][00];
		//diff_pixel[02][00][01] <= numero[00][01] > 58 ? numero[00][01] - 58 : 58 - numero[00][01];
		//diff_pixel[02][00][02] <= numero[00][02] > 80 ? numero[00][02] - 80 : 80 - numero[00][02];
		//diff_pixel[02][00][03] <= numero[00][03] > 101 ? numero[00][03] - 101 : 101 - numero[00][03];
		//diff_pixel[02][00][04] <= numero[00][04] > 101 ? numero[00][04] - 101 : 101 - numero[00][04];
		//diff_pixel[02][00][05] <= numero[00][05] > 103 ? numero[00][05] - 103 : 103 - numero[00][05];
		//diff_pixel[02][00][06] <= numero[00][06] > 99 ? numero[00][06] - 99 : 99 - numero[00][06];
		//diff_pixel[02][00][07] <= numero[00][07] > 92 ? numero[00][07] - 92 : 92 - numero[00][07];
		//diff_pixel[02][00][08] <= numero[00][08] > 76 ? numero[00][08] - 76 : 76 - numero[00][08];
		//diff_pixel[02][00][09] <= numero[00][09] > 51 ? numero[00][09] - 51 : 51 - numero[00][09];
		//diff_pixel[02][00][10] <= numero[00][10] > 22 ? numero[00][10] - 22 : 22 - numero[00][10];
		//diff_pixel[02][01][00] <= numero[01][00] > 46 ? numero[01][00] - 46 : 46 - numero[01][00];
		//diff_pixel[02][01][01] <= numero[01][01] > 89 ? numero[01][01] - 89 : 89 - numero[01][01];
		//diff_pixel[02][01][02] <= numero[01][02] > 126 ? numero[01][02] - 126 : 126 - numero[01][02];
		//diff_pixel[02][01][03] <= numero[01][03] > 143 ? numero[01][03] - 143 : 143 - numero[01][03];
		//diff_pixel[02][01][04] <= numero[01][04] > 143 ? numero[01][04] - 143 : 143 - numero[01][04];
		//diff_pixel[02][01][05] <= numero[01][05] > 138 ? numero[01][05] - 138 : 138 - numero[01][05];
		//diff_pixel[02][01][06] <= numero[01][06] > 142 ? numero[01][06] - 142 : 142 - numero[01][06];
		//diff_pixel[02][01][07] <= numero[01][07] > 140 ? numero[01][07] - 140 : 140 - numero[01][07];
		//diff_pixel[02][01][08] <= numero[01][08] > 135 ? numero[01][08] - 135 : 135 - numero[01][08];
		//diff_pixel[02][01][09] <= numero[01][09] > 107 ? numero[01][09] - 107 : 107 - numero[01][09];
		//diff_pixel[02][01][10] <= numero[01][10] > 62 ? numero[01][10] - 62 : 62 - numero[01][10];
		diff_pixel[02][02][00] <= numero[02][00] > 98 ? numero[02][00] - 98 : 98 - numero[02][00];
		diff_pixel[02][02][01] <= numero[02][01] > 123 ? numero[02][01] - 123 : 123 - numero[02][01];
		diff_pixel[02][02][02] <= numero[02][02] > 117 ? numero[02][02] - 117 : 117 - numero[02][02];
		diff_pixel[02][02][03] <= numero[02][03] > 80 ? numero[02][03] - 80 : 80 - numero[02][03];
		diff_pixel[02][02][04] <= numero[02][04] > 31 ? numero[02][04] - 31 : 31 - numero[02][04];
		diff_pixel[02][02][05] <= numero[02][05] > 9 ? numero[02][05] - 9 : 9 - numero[02][05];
		diff_pixel[02][02][06] <= numero[02][06] > 23 ? numero[02][06] - 23 : 23 - numero[02][06];
		diff_pixel[02][02][07] <= numero[02][07] > 60 ? numero[02][07] - 60 : 60 - numero[02][07];
		diff_pixel[02][02][08] <= numero[02][08] > 107 ? numero[02][08] - 107 : 107 - numero[02][08];
		diff_pixel[02][02][09] <= numero[02][09] > 125 ? numero[02][09] - 125 : 125 - numero[02][09];
		diff_pixel[02][02][10] <= numero[02][10] > 114 ? numero[02][10] - 114 : 114 - numero[02][10];
		diff_pixel[02][03][00] <= numero[03][00] > 31 ? numero[03][00] - 31 : 31 - numero[03][00];
		diff_pixel[02][03][01] <= numero[03][01] > 43 ? numero[03][01] - 43 : 43 - numero[03][01];
		diff_pixel[02][03][02] <= numero[03][02] > 38 ? numero[03][02] - 38 : 38 - numero[03][02];
		diff_pixel[02][03][03] <= numero[03][03] > 21 ? numero[03][03] - 21 : 21 - numero[03][03];
		diff_pixel[02][03][04] <= numero[03][04] > 9 ? numero[03][04] - 9 : 9 - numero[03][04];
		diff_pixel[02][03][05] <= numero[03][05] > 18 ? numero[03][05] - 18 : 18 - numero[03][05];
		diff_pixel[02][03][06] <= numero[03][06] > 54 ? numero[03][06] - 54 : 54 - numero[03][06];
		diff_pixel[02][03][07] <= numero[03][07] > 101 ? numero[03][07] - 101 : 101 - numero[03][07];
		diff_pixel[02][03][08] <= numero[03][08] > 141 ? numero[03][08] - 141 : 141 - numero[03][08];
		diff_pixel[02][03][09] <= numero[03][09] > 142 ? numero[03][09] - 142 : 142 - numero[03][09];
		diff_pixel[02][03][10] <= numero[03][10] > 126 ? numero[03][10] - 126 : 126 - numero[03][10];
		diff_pixel[02][04][00] <= numero[04][00] > 0 ? numero[04][00] - 0 : 0 - numero[04][00];
		diff_pixel[02][04][01] <= numero[04][01] > 0 ? numero[04][01] - 0 : 0 - numero[04][01];
		diff_pixel[02][04][02] <= numero[04][02] > 6 ? numero[04][02] - 6 : 6 - numero[04][02];
		diff_pixel[02][04][03] <= numero[04][03] > 22 ? numero[04][03] - 22 : 22 - numero[04][03];
		diff_pixel[02][04][04] <= numero[04][04] > 48 ? numero[04][04] - 48 : 48 - numero[04][04];
		diff_pixel[02][04][05] <= numero[04][05] > 76 ? numero[04][05] - 76 : 76 - numero[04][05];
		diff_pixel[02][04][06] <= numero[04][06] > 116 ? numero[04][06] - 116 : 116 - numero[04][06];
		diff_pixel[02][04][07] <= numero[04][07] > 146 ? numero[04][07] - 146 : 146 - numero[04][07];
		diff_pixel[02][04][08] <= numero[04][08] > 160 ? numero[04][08] - 160 : 160 - numero[04][08];
		diff_pixel[02][04][09] <= numero[04][09] > 139 ? numero[04][09] - 139 : 139 - numero[04][09];
		diff_pixel[02][04][10] <= numero[04][10] > 114 ? numero[04][10] - 114 : 114 - numero[04][10];
		diff_pixel[02][05][00] <= numero[05][00] > 8 ? numero[05][00] - 8 : 8 - numero[05][00];
		diff_pixel[02][05][01] <= numero[05][01] > 10 ? numero[05][01] - 10 : 10 - numero[05][01];
		diff_pixel[02][05][02] <= numero[05][02] > 39 ? numero[05][02] - 39 : 39 - numero[05][02];
		diff_pixel[02][05][03] <= numero[05][03] > 89 ? numero[05][03] - 89 : 89 - numero[05][03];
		diff_pixel[02][05][04] <= numero[05][04] > 133 ? numero[05][04] - 133 : 133 - numero[05][04];
		diff_pixel[02][05][05] <= numero[05][05] > 159 ? numero[05][05] - 159 : 159 - numero[05][05];
		diff_pixel[02][05][06] <= numero[05][06] > 179 ? numero[05][06] - 179 : 179 - numero[05][06];
		diff_pixel[02][05][07] <= numero[05][07] > 169 ? numero[05][07] - 169 : 169 - numero[05][07];
		diff_pixel[02][05][08] <= numero[05][08] > 145 ? numero[05][08] - 145 : 145 - numero[05][08];
		diff_pixel[02][05][09] <= numero[05][09] > 102 ? numero[05][09] - 102 : 102 - numero[05][09];
		diff_pixel[02][05][10] <= numero[05][10] > 63 ? numero[05][10] - 63 : 63 - numero[05][10];
		diff_pixel[02][06][00] <= numero[06][00] > 26 ? numero[06][00] - 26 : 26 - numero[06][00];
		diff_pixel[02][06][01] <= numero[06][01] > 44 ? numero[06][01] - 44 : 44 - numero[06][01];
		diff_pixel[02][06][02] <= numero[06][02] > 92 ? numero[06][02] - 92 : 92 - numero[06][02];
		diff_pixel[02][06][03] <= numero[06][03] > 138 ? numero[06][03] - 138 : 138 - numero[06][03];
		diff_pixel[02][06][04] <= numero[06][04] > 170 ? numero[06][04] - 170 : 170 - numero[06][04];
		diff_pixel[02][06][05] <= numero[06][05] > 177 ? numero[06][05] - 177 : 177 - numero[06][05];
		diff_pixel[02][06][06] <= numero[06][06] > 167 ? numero[06][06] - 167 : 167 - numero[06][06];
		diff_pixel[02][06][07] <= numero[06][07] > 138 ? numero[06][07] - 138 : 138 - numero[06][07];
		diff_pixel[02][06][08] <= numero[06][08] > 93 ? numero[06][08] - 93 : 93 - numero[06][08];
		diff_pixel[02][06][09] <= numero[06][09] > 50 ? numero[06][09] - 50 : 50 - numero[06][09];
		diff_pixel[02][06][10] <= numero[06][10] > 24 ? numero[06][10] - 24 : 24 - numero[06][10];
		diff_pixel[02][07][00] <= numero[07][00] > 62 ? numero[07][00] - 62 : 62 - numero[07][00];
		diff_pixel[02][07][01] <= numero[07][01] > 89 ? numero[07][01] - 89 : 89 - numero[07][01];
		diff_pixel[02][07][02] <= numero[07][02] > 132 ? numero[07][02] - 132 : 132 - numero[07][02];
		diff_pixel[02][07][03] <= numero[07][03] > 156 ? numero[07][03] - 156 : 156 - numero[07][03];
		diff_pixel[02][07][04] <= numero[07][04] > 159 ? numero[07][04] - 159 : 159 - numero[07][04];
		diff_pixel[02][07][05] <= numero[07][05] > 139 ? numero[07][05] - 139 : 139 - numero[07][05];
		diff_pixel[02][07][06] <= numero[07][06] > 111 ? numero[07][06] - 111 : 111 - numero[07][06];
		diff_pixel[02][07][07] <= numero[07][07] > 79 ? numero[07][07] - 79 : 79 - numero[07][07];
		diff_pixel[02][07][08] <= numero[07][08] > 44 ? numero[07][08] - 44 : 44 - numero[07][08];
		diff_pixel[02][07][09] <= numero[07][09] > 15 ? numero[07][09] - 15 : 15 - numero[07][09];
		diff_pixel[02][07][10] <= numero[07][10] > 5 ? numero[07][10] - 5 : 5 - numero[07][10];
		//diff_pixel[02][08][00] <= numero[08][00] > 123 ? numero[08][00] - 123 : 123 - numero[08][00];
		//diff_pixel[02][08][01] <= numero[08][01] > 151 ? numero[08][01] - 151 : 151 - numero[08][01];
		//diff_pixel[02][08][02] <= numero[08][02] > 166 ? numero[08][02] - 166 : 166 - numero[08][02];
		//diff_pixel[02][08][03] <= numero[08][03] > 153 ? numero[08][03] - 153 : 153 - numero[08][03];
		//diff_pixel[02][08][04] <= numero[08][04] > 109 ? numero[08][04] - 109 : 109 - numero[08][04];
		//diff_pixel[02][08][05] <= numero[08][05] > 52 ? numero[08][05] - 52 : 52 - numero[08][05];
		//diff_pixel[02][08][06] <= numero[08][06] > 11 ? numero[08][06] - 11 : 11 - numero[08][06];
		//diff_pixel[02][08][07] <= numero[08][07] > 0 ? numero[08][07] - 0 : 0 - numero[08][07];
		//diff_pixel[02][08][08] <= numero[08][08] > 0 ? numero[08][08] - 0 : 0 - numero[08][08];
		//diff_pixel[02][08][09] <= numero[08][09] > 0 ? numero[08][09] - 0 : 0 - numero[08][09];
		//diff_pixel[02][08][10] <= numero[08][10] > 0 ? numero[08][10] - 0 : 0 - numero[08][10];
		//diff_pixel[02][09][00] <= numero[09][00] > 106 ? numero[09][00] - 106 : 106 - numero[09][00];
		//diff_pixel[02][09][01] <= numero[09][01] > 149 ? numero[09][01] - 149 : 149 - numero[09][01];
		//diff_pixel[02][09][02] <= numero[09][02] > 173 ? numero[09][02] - 173 : 173 - numero[09][02];
		//diff_pixel[02][09][03] <= numero[09][03] > 175 ? numero[09][03] - 175 : 175 - numero[09][03];
		//diff_pixel[02][09][04] <= numero[09][04] > 161 ? numero[09][04] - 161 : 161 - numero[09][04];
		//diff_pixel[02][09][05] <= numero[09][05] > 142 ? numero[09][05] - 142 : 142 - numero[09][05];
		//diff_pixel[02][09][06] <= numero[09][06] > 129 ? numero[09][06] - 129 : 129 - numero[09][06];
		//diff_pixel[02][09][07] <= numero[09][07] > 123 ? numero[09][07] - 123 : 123 - numero[09][07];
		//diff_pixel[02][09][08] <= numero[09][08] > 118 ? numero[09][08] - 118 : 118 - numero[09][08];
		//diff_pixel[02][09][09] <= numero[09][09] > 104 ? numero[09][09] - 104 : 104 - numero[09][09];
		//diff_pixel[02][09][10] <= numero[09][10] > 79 ? numero[09][10] - 79 : 79 - numero[09][10];
		//diff_pixel[02][10][00] <= numero[10][00] > 68 ? numero[10][00] - 68 : 68 - numero[10][00];
		//diff_pixel[02][10][01] <= numero[10][01] > 103 ? numero[10][01] - 103 : 103 - numero[10][01];
		//diff_pixel[02][10][02] <= numero[10][02] > 118 ? numero[10][02] - 118 : 118 - numero[10][02];
		//diff_pixel[02][10][03] <= numero[10][03] > 125 ? numero[10][03] - 125 : 125 - numero[10][03];
		//diff_pixel[02][10][04] <= numero[10][04] > 121 ? numero[10][04] - 121 : 121 - numero[10][04];
		//diff_pixel[02][10][05] <= numero[10][05] > 120 ? numero[10][05] - 120 : 120 - numero[10][05];
		//diff_pixel[02][10][06] <= numero[10][06] > 120 ? numero[10][06] - 120 : 120 - numero[10][06];
		//diff_pixel[02][10][07] <= numero[10][07] > 121 ? numero[10][07] - 121 : 121 - numero[10][07];
		//diff_pixel[02][10][08] <= numero[10][08] > 116 ? numero[10][08] - 116 : 116 - numero[10][08];
		//diff_pixel[02][10][09] <= numero[10][09] > 100 ? numero[10][09] - 100 : 100 - numero[10][09];
		//diff_pixel[02][10][10] <= numero[10][10] > 80 ? numero[10][10] - 80 : 80 - numero[10][10];
		
		//diff_pixel[03][00][00] <= numero[00][00] > 24 ? numero[00][00] - 24 : 24 - numero[00][00];
		//diff_pixel[03][00][01] <= numero[00][01] > 39 ? numero[00][01] - 39 : 39 - numero[00][01];
		//diff_pixel[03][00][02] <= numero[00][02] > 67 ? numero[00][02] - 67 : 67 - numero[00][02];
		//diff_pixel[03][00][03] <= numero[00][03] > 90 ? numero[00][03] - 90 : 90 - numero[00][03];
		//diff_pixel[03][00][04] <= numero[00][04] > 98 ? numero[00][04] - 98 : 98 - numero[00][04];
		//diff_pixel[03][00][05] <= numero[00][05] > 100 ? numero[00][05] - 100 : 100 - numero[00][05];
		//diff_pixel[03][00][06] <= numero[00][06] > 98 ? numero[00][06] - 98 : 98 - numero[00][06];
		//diff_pixel[03][00][07] <= numero[00][07] > 98 ? numero[00][07] - 98 : 98 - numero[00][07];
		//diff_pixel[03][00][08] <= numero[00][08] > 96 ? numero[00][08] - 96 : 96 - numero[00][08];
		//diff_pixel[03][00][09] <= numero[00][09] > 83 ? numero[00][09] - 83 : 83 - numero[00][09];
		//diff_pixel[03][00][10] <= numero[00][10] > 64 ? numero[00][10] - 64 : 64 - numero[00][10];
		//diff_pixel[03][01][00] <= numero[01][00] > 32 ? numero[01][00] - 32 : 32 - numero[01][00];
		//diff_pixel[03][01][01] <= numero[01][01] > 54 ? numero[01][01] - 54 : 54 - numero[01][01];
		//diff_pixel[03][01][02] <= numero[01][02] > 91 ? numero[01][02] - 91 : 91 - numero[01][02];
		//diff_pixel[03][01][03] <= numero[01][03] > 121 ? numero[01][03] - 121 : 121 - numero[01][03];
		//diff_pixel[03][01][04] <= numero[01][04] > 138 ? numero[01][04] - 138 : 138 - numero[01][04];
		//diff_pixel[03][01][05] <= numero[01][05] > 146 ? numero[01][05] - 146 : 146 - numero[01][05];
		//diff_pixel[03][01][06] <= numero[01][06] > 157 ? numero[01][06] - 157 : 157 - numero[01][06];
		//diff_pixel[03][01][07] <= numero[01][07] > 166 ? numero[01][07] - 166 : 166 - numero[01][07];
		//diff_pixel[03][01][08] <= numero[01][08] > 164 ? numero[01][08] - 164 : 164 - numero[01][08];
		//diff_pixel[03][01][09] <= numero[01][09] > 139 ? numero[01][09] - 139 : 139 - numero[01][09];
		//diff_pixel[03][01][10] <= numero[01][10] > 99 ? numero[01][10] - 99 : 99 - numero[01][10];
		diff_pixel[03][02][00] <= numero[02][00] > 0 ? numero[02][00] - 0 : 0 - numero[02][00];
		diff_pixel[03][02][01] <= numero[02][01] > 1 ? numero[02][01] - 1 : 1 - numero[02][01];
		diff_pixel[03][02][02] <= numero[02][02] > 5 ? numero[02][02] - 5 : 5 - numero[02][02];
		diff_pixel[03][02][03] <= numero[02][03] > 6 ? numero[02][03] - 6 : 6 - numero[02][03];
		diff_pixel[03][02][04] <= numero[02][04] > 21 ? numero[02][04] - 21 : 21 - numero[02][04];
		diff_pixel[03][02][05] <= numero[02][05] > 48 ? numero[02][05] - 48 : 48 - numero[02][05];
		diff_pixel[03][02][06] <= numero[02][06] > 94 ? numero[02][06] - 94 : 94 - numero[02][06];
		diff_pixel[03][02][07] <= numero[02][07] > 127 ? numero[02][07] - 127 : 127 - numero[02][07];
		diff_pixel[03][02][08] <= numero[02][08] > 130 ? numero[02][08] - 130 : 130 - numero[02][08];
		diff_pixel[03][02][09] <= numero[02][09] > 102 ? numero[02][09] - 102 : 102 - numero[02][09];
		diff_pixel[03][02][10] <= numero[02][10] > 51 ? numero[02][10] - 51 : 51 - numero[02][10];
		diff_pixel[03][03][00] <= numero[03][00] > 0 ? numero[03][00] - 0 : 0 - numero[03][00];
		diff_pixel[03][03][01] <= numero[03][01] > 0 ? numero[03][01] - 0 : 0 - numero[03][01];
		diff_pixel[03][03][02] <= numero[03][02] > 0 ? numero[03][02] - 0 : 0 - numero[03][02];
		diff_pixel[03][03][03] <= numero[03][03] > 13 ? numero[03][03] - 13 : 13 - numero[03][03];
		diff_pixel[03][03][04] <= numero[03][04] > 43 ? numero[03][04] - 43 : 43 - numero[03][04];
		diff_pixel[03][03][05] <= numero[03][05] > 83 ? numero[03][05] - 83 : 83 - numero[03][05];
		diff_pixel[03][03][06] <= numero[03][06] > 113 ? numero[03][06] - 113 : 113 - numero[03][06];
		diff_pixel[03][03][07] <= numero[03][07] > 115 ? numero[03][07] - 115 : 115 - numero[03][07];
		diff_pixel[03][03][08] <= numero[03][08] > 88 ? numero[03][08] - 88 : 88 - numero[03][08];
		diff_pixel[03][03][09] <= numero[03][09] > 48 ? numero[03][09] - 48 : 48 - numero[03][09];
		diff_pixel[03][03][10] <= numero[03][10] > 22 ? numero[03][10] - 22 : 22 - numero[03][10];
		diff_pixel[03][04][00] <= numero[04][00] > 0 ? numero[04][00] - 0 : 0 - numero[04][00];
		diff_pixel[03][04][01] <= numero[04][01] > 0 ? numero[04][01] - 0 : 0 - numero[04][01];
		diff_pixel[03][04][02] <= numero[04][02] > 19 ? numero[04][02] - 19 : 19 - numero[04][02];
		diff_pixel[03][04][03] <= numero[04][03] > 53 ? numero[04][03] - 53 : 53 - numero[04][03];
		diff_pixel[03][04][04] <= numero[04][04] > 94 ? numero[04][04] - 94 : 94 - numero[04][04];
		diff_pixel[03][04][05] <= numero[04][05] > 136 ? numero[04][05] - 136 : 136 - numero[04][05];
		diff_pixel[03][04][06] <= numero[04][06] > 149 ? numero[04][06] - 149 : 149 - numero[04][06];
		diff_pixel[03][04][07] <= numero[04][07] > 133 ? numero[04][07] - 133 : 133 - numero[04][07];
		diff_pixel[03][04][08] <= numero[04][08] > 88 ? numero[04][08] - 88 : 88 - numero[04][08];
		diff_pixel[03][04][09] <= numero[04][09] > 42 ? numero[04][09] - 42 : 42 - numero[04][09];
		diff_pixel[03][04][10] <= numero[04][10] > 21 ? numero[04][10] - 21 : 21 - numero[04][10];
		diff_pixel[03][05][00] <= numero[05][00] > 0 ? numero[05][00] - 0 : 0 - numero[05][00];
		diff_pixel[03][05][01] <= numero[05][01] > 12 ? numero[05][01] - 12 : 12 - numero[05][01];
		diff_pixel[03][05][02] <= numero[05][02] > 45 ? numero[05][02] - 45 : 45 - numero[05][02];
		diff_pixel[03][05][03] <= numero[05][03] > 94 ? numero[05][03] - 94 : 94 - numero[05][03];
		diff_pixel[03][05][04] <= numero[05][04] > 138 ? numero[05][04] - 138 : 138 - numero[05][04];
		diff_pixel[03][05][05] <= numero[05][05] > 166 ? numero[05][05] - 166 : 166 - numero[05][05];
		diff_pixel[03][05][06] <= numero[05][06] > 184 ? numero[05][06] - 184 : 184 - numero[05][06];
		diff_pixel[03][05][07] <= numero[05][07] > 169 ? numero[05][07] - 169 : 169 - numero[05][07];
		diff_pixel[03][05][08] <= numero[05][08] > 142 ? numero[05][08] - 142 : 142 - numero[05][08];
		diff_pixel[03][05][09] <= numero[05][09] > 96 ? numero[05][09] - 96 : 96 - numero[05][09];
		diff_pixel[03][05][10] <= numero[05][10] > 57 ? numero[05][10] - 57 : 57 - numero[05][10];
		diff_pixel[03][06][00] <= numero[06][00] > 2 ? numero[06][00] - 2 : 2 - numero[06][00];
		diff_pixel[03][06][01] <= numero[06][01] > 0 ? numero[06][01] - 0 : 0 - numero[06][01];
		diff_pixel[03][06][02] <= numero[06][02] > 12 ? numero[06][02] - 12 : 12 - numero[06][02];
		diff_pixel[03][06][03] <= numero[06][03] > 32 ? numero[06][03] - 32 : 32 - numero[06][03];
		diff_pixel[03][06][04] <= numero[06][04] > 49 ? numero[06][04] - 49 : 49 - numero[06][04];
		diff_pixel[03][06][05] <= numero[06][05] > 61 ? numero[06][05] - 61 : 61 - numero[06][05];
		diff_pixel[03][06][06] <= numero[06][06] > 81 ? numero[06][06] - 81 : 81 - numero[06][06];
		diff_pixel[03][06][07] <= numero[06][07] > 99 ? numero[06][07] - 99 : 99 - numero[06][07];
		diff_pixel[03][06][08] <= numero[06][08] > 117 ? numero[06][08] - 117 : 117 - numero[06][08];
		diff_pixel[03][06][09] <= numero[06][09] > 110 ? numero[06][09] - 110 : 110 - numero[06][09];
		diff_pixel[03][06][10] <= numero[06][10] > 99 ? numero[06][10] - 99 : 99 - numero[06][10];
		diff_pixel[03][07][00] <= numero[07][00] > 38 ? numero[07][00] - 38 : 38 - numero[07][00];
		diff_pixel[03][07][01] <= numero[07][01] > 26 ? numero[07][01] - 26 : 26 - numero[07][01];
		diff_pixel[03][07][02] <= numero[07][02] > 23 ? numero[07][02] - 23 : 23 - numero[07][02];
		diff_pixel[03][07][03] <= numero[07][03] > 14 ? numero[07][03] - 14 : 14 - numero[07][03];
		diff_pixel[03][07][04] <= numero[07][04] > 0 ? numero[07][04] - 0 : 0 - numero[07][04];
		diff_pixel[03][07][05] <= numero[07][05] > 0 ? numero[07][05] - 0 : 0 - numero[07][05];
		diff_pixel[03][07][06] <= numero[07][06] > 22 ? numero[07][06] - 22 : 22 - numero[07][06];
		diff_pixel[03][07][07] <= numero[07][07] > 59 ? numero[07][07] - 59 : 59 - numero[07][07];
		diff_pixel[03][07][08] <= numero[07][08] > 110 ? numero[07][08] - 110 : 110 - numero[07][08];
		diff_pixel[03][07][09] <= numero[07][09] > 126 ? numero[07][09] - 126 : 126 - numero[07][09];
		diff_pixel[03][07][10] <= numero[07][10] > 125 ? numero[07][10] - 125 : 125 - numero[07][10];
		//diff_pixel[03][08][00] <= numero[08][00] > 129 ? numero[08][00] - 129 : 129 - numero[08][00];
		//diff_pixel[03][08][01] <= numero[08][01] > 131 ? numero[08][01] - 131 : 131 - numero[08][01];
		//diff_pixel[03][08][02] <= numero[08][02] > 119 ? numero[08][02] - 119 : 119 - numero[08][02];
		//diff_pixel[03][08][03] <= numero[08][03] > 80 ? numero[08][03] - 80 : 80 - numero[08][03];
		//diff_pixel[03][08][04] <= numero[08][04] > 30 ? numero[08][04] - 30 : 30 - numero[08][04];
		//diff_pixel[03][08][05] <= numero[08][05] > 6 ? numero[08][05] - 6 : 6 - numero[08][05];
		//diff_pixel[03][08][06] <= numero[08][06] > 16 ? numero[08][06] - 16 : 16 - numero[08][06];
		//diff_pixel[03][08][07] <= numero[08][07] > 56 ? numero[08][07] - 56 : 56 - numero[08][07];
		//diff_pixel[03][08][08] <= numero[08][08] > 102 ? numero[08][08] - 102 : 102 - numero[08][08];
		//diff_pixel[03][08][09] <= numero[08][09] > 119 ? numero[08][09] - 119 : 119 - numero[08][09];
		//diff_pixel[03][08][10] <= numero[08][10] > 110 ? numero[08][10] - 110 : 110 - numero[08][10];
		//diff_pixel[03][09][00] <= numero[09][00] > 54 ? numero[09][00] - 54 : 54 - numero[09][00];
		//diff_pixel[03][09][01] <= numero[09][01] > 88 ? numero[09][01] - 88 : 88 - numero[09][01];
		//diff_pixel[03][09][02] <= numero[09][02] > 120 ? numero[09][02] - 120 : 120 - numero[09][02];
		//diff_pixel[03][09][03] <= numero[09][03] > 132 ? numero[09][03] - 132 : 132 - numero[09][03];
		//diff_pixel[03][09][04] <= numero[09][04] > 127 ? numero[09][04] - 127 : 127 - numero[09][04];
		//diff_pixel[03][09][05] <= numero[09][05] > 122 ? numero[09][05] - 122 : 122 - numero[09][05];
		//diff_pixel[03][09][06] <= numero[09][06] > 124 ? numero[09][06] - 124 : 124 - numero[09][06];
		//diff_pixel[03][09][07] <= numero[09][07] > 126 ? numero[09][07] - 126 : 126 - numero[09][07];
		//diff_pixel[03][09][08] <= numero[09][08] > 125 ? numero[09][08] - 125 : 125 - numero[09][08];
		//diff_pixel[03][09][09] <= numero[09][09] > 99 ? numero[09][09] - 99 : 99 - numero[09][09];
		//diff_pixel[03][09][10] <= numero[09][10] > 65 ? numero[09][10] - 65 : 65 - numero[09][10];
		//diff_pixel[03][10][00] <= numero[10][00] > 23 ? numero[10][00] - 23 : 23 - numero[10][00];
		//diff_pixel[03][10][01] <= numero[10][01] > 56 ? numero[10][01] - 56 : 56 - numero[10][01];
		//diff_pixel[03][10][02] <= numero[10][02] > 92 ? numero[10][02] - 92 : 92 - numero[10][02];
		//diff_pixel[03][10][03] <= numero[10][03] > 116 ? numero[10][03] - 116 : 116 - numero[10][03];
		//diff_pixel[03][10][04] <= numero[10][04] > 128 ? numero[10][04] - 128 : 128 - numero[10][04];
		//diff_pixel[03][10][05] <= numero[10][05] > 130 ? numero[10][05] - 130 : 130 - numero[10][05];
		//diff_pixel[03][10][06] <= numero[10][06] > 126 ? numero[10][06] - 126 : 126 - numero[10][06];
		//diff_pixel[03][10][07] <= numero[10][07] > 115 ? numero[10][07] - 115 : 115 - numero[10][07];
		//diff_pixel[03][10][08] <= numero[10][08] > 94 ? numero[10][08] - 94 : 94 - numero[10][08];
		//diff_pixel[03][10][09] <= numero[10][09] > 63 ? numero[10][09] - 63 : 63 - numero[10][09];
		//diff_pixel[03][10][10] <= numero[10][10] > 24 ? numero[10][10] - 24 : 24 - numero[10][10];
		
		//diff_pixel[04][00][00] <= numero[00][00] > 14 ? numero[00][00] - 14 : 14 - numero[00][00];
		//diff_pixel[04][00][01] <= numero[00][01] > 14 ? numero[00][01] - 14 : 14 - numero[00][01];
		//diff_pixel[04][00][02] <= numero[00][02] > 10 ? numero[00][02] - 10 : 10 - numero[00][02];
		//diff_pixel[04][00][03] <= numero[00][03] > 24 ? numero[00][03] - 24 : 24 - numero[00][03];
		//diff_pixel[04][00][04] <= numero[00][04] > 40 ? numero[00][04] - 40 : 40 - numero[00][04];
		//diff_pixel[04][00][05] <= numero[00][05] > 70 ? numero[00][05] - 70 : 70 - numero[00][05];
		//diff_pixel[04][00][06] <= numero[00][06] > 89 ? numero[00][06] - 89 : 89 - numero[00][06];
		//diff_pixel[04][00][07] <= numero[00][07] > 91 ? numero[00][07] - 91 : 91 - numero[00][07];
		//diff_pixel[04][00][08] <= numero[00][08] > 78 ? numero[00][08] - 78 : 78 - numero[00][08];
		//diff_pixel[04][00][09] <= numero[00][09] > 50 ? numero[00][09] - 50 : 50 - numero[00][09];
		//diff_pixel[04][00][10] <= numero[00][10] > 19 ? numero[00][10] - 19 : 19 - numero[00][10];
		//diff_pixel[04][01][00] <= numero[01][00] > 0 ? numero[01][00] - 0 : 0 - numero[01][00];
		//diff_pixel[04][01][01] <= numero[01][01] > 0 ? numero[01][01] - 0 : 0 - numero[01][01];
		//diff_pixel[04][01][02] <= numero[01][02] > 12 ? numero[01][02] - 12 : 12 - numero[01][02];
		//diff_pixel[04][01][03] <= numero[01][03] > 46 ? numero[01][03] - 46 : 46 - numero[01][03];
		//diff_pixel[04][01][04] <= numero[01][04] > 86 ? numero[01][04] - 86 : 86 - numero[01][04];
		//diff_pixel[04][01][05] <= numero[01][05] > 134 ? numero[01][05] - 134 : 134 - numero[01][05];
		//diff_pixel[04][01][06] <= numero[01][06] > 166 ? numero[01][06] - 166 : 166 - numero[01][06];
		//diff_pixel[04][01][07] <= numero[01][07] > 167 ? numero[01][07] - 167 : 167 - numero[01][07];
		//diff_pixel[04][01][08] <= numero[01][08] > 143 ? numero[01][08] - 143 : 143 - numero[01][08];
		//diff_pixel[04][01][09] <= numero[01][09] > 95 ? numero[01][09] - 95 : 95 - numero[01][09];
		//diff_pixel[04][01][10] <= numero[01][10] > 44 ? numero[01][10] - 44 : 44 - numero[01][10];
		diff_pixel[04][02][00] <= numero[02][00] > 0 ? numero[02][00] - 0 : 0 - numero[02][00];
		diff_pixel[04][02][01] <= numero[02][01] > 20 ? numero[02][01] - 20 : 20 - numero[02][01];
		diff_pixel[04][02][02] <= numero[02][02] > 49 ? numero[02][02] - 49 : 49 - numero[02][02];
		diff_pixel[04][02][03] <= numero[02][03] > 98 ? numero[02][03] - 98 : 98 - numero[02][03];
		diff_pixel[04][02][04] <= numero[02][04] > 139 ? numero[02][04] - 139 : 139 - numero[02][04];
		diff_pixel[04][02][05] <= numero[02][05] > 168 ? numero[02][05] - 168 : 168 - numero[02][05];
		diff_pixel[04][02][06] <= numero[02][06] > 182 ? numero[02][06] - 182 : 182 - numero[02][06];
		diff_pixel[04][02][07] <= numero[02][07] > 168 ? numero[02][07] - 168 : 168 - numero[02][07];
		diff_pixel[04][02][08] <= numero[02][08] > 136 ? numero[02][08] - 136 : 136 - numero[02][08];
		diff_pixel[04][02][09] <= numero[02][09] > 91 ? numero[02][09] - 91 : 91 - numero[02][09];
		diff_pixel[04][02][10] <= numero[02][10] > 44 ? numero[02][10] - 44 : 44 - numero[02][10];
		diff_pixel[04][03][00] <= numero[03][00] > 24 ? numero[03][00] - 24 : 24 - numero[03][00];
		diff_pixel[04][03][01] <= numero[03][01] > 51 ? numero[03][01] - 51 : 51 - numero[03][01];
		diff_pixel[04][03][02] <= numero[03][02] > 91 ? numero[03][02] - 91 : 91 - numero[03][02];
		diff_pixel[04][03][03] <= numero[03][03] > 117 ? numero[03][03] - 117 : 117 - numero[03][03];
		diff_pixel[04][03][04] <= numero[03][04] > 132 ? numero[03][04] - 132 : 132 - numero[03][04];
		diff_pixel[04][03][05] <= numero[03][05] > 127 ? numero[03][05] - 127 : 127 - numero[03][05];
		diff_pixel[04][03][06] <= numero[03][06] > 136 ? numero[03][06] - 136 : 136 - numero[03][06];
		diff_pixel[04][03][07] <= numero[03][07] > 139 ? numero[03][07] - 139 : 139 - numero[03][07];
		diff_pixel[04][03][08] <= numero[03][08] > 126 ? numero[03][08] - 126 : 126 - numero[03][08];
		diff_pixel[04][03][09] <= numero[03][09] > 93 ? numero[03][09] - 93 : 93 - numero[03][09];
		diff_pixel[04][03][10] <= numero[03][10] > 51 ? numero[03][10] - 51 : 51 - numero[03][10];
		diff_pixel[04][04][00] <= numero[04][00] > 78 ? numero[04][00] - 78 : 78 - numero[04][00];
		diff_pixel[04][04][01] <= numero[04][01] > 98 ? numero[04][01] - 98 : 98 - numero[04][01];
		diff_pixel[04][04][02] <= numero[04][02] > 116 ? numero[04][02] - 116 : 116 - numero[04][02];
		diff_pixel[04][04][03] <= numero[04][03] > 112 ? numero[04][03] - 112 : 112 - numero[04][03];
		diff_pixel[04][04][04] <= numero[04][04] > 92 ? numero[04][04] - 92 : 92 - numero[04][04];
		diff_pixel[04][04][05] <= numero[04][05] > 77 ? numero[04][05] - 77 : 77 - numero[04][05];
		diff_pixel[04][04][06] <= numero[04][06] > 99 ? numero[04][06] - 99 : 99 - numero[04][06];
		diff_pixel[04][04][07] <= numero[04][07] > 120 ? numero[04][07] - 120 : 120 - numero[04][07];
		diff_pixel[04][04][08] <= numero[04][08] > 126 ? numero[04][08] - 126 : 126 - numero[04][08];
		diff_pixel[04][04][09] <= numero[04][09] > 97 ? numero[04][09] - 97 : 97 - numero[04][09];
		diff_pixel[04][04][10] <= numero[04][10] > 63 ? numero[04][10] - 63 : 63 - numero[04][10];
		diff_pixel[04][05][00] <= numero[05][00] > 123 ? numero[05][00] - 123 : 123 - numero[05][00];
		diff_pixel[04][05][01] <= numero[05][01] > 128 ? numero[05][01] - 128 : 128 - numero[05][01];
		diff_pixel[04][05][02] <= numero[05][02] > 119 ? numero[05][02] - 119 : 119 - numero[05][02];
		diff_pixel[04][05][03] <= numero[05][03] > 84 ? numero[05][03] - 84 : 84 - numero[05][03];
		diff_pixel[04][05][04] <= numero[05][04] > 52 ? numero[05][04] - 52 : 52 - numero[05][04];
		diff_pixel[04][05][05] <= numero[05][05] > 51 ? numero[05][05] - 51 : 51 - numero[05][05];
		diff_pixel[04][05][06] <= numero[05][06] > 86 ? numero[05][06] - 86 : 86 - numero[05][06];
		diff_pixel[04][05][07] <= numero[05][07] > 123 ? numero[05][07] - 123 : 123 - numero[05][07];
		diff_pixel[04][05][08] <= numero[05][08] > 128 ? numero[05][08] - 128 : 128 - numero[05][08];
		diff_pixel[04][05][09] <= numero[05][09] > 97 ? numero[05][09] - 97 : 97 - numero[05][09];
		diff_pixel[04][05][10] <= numero[05][10] > 59 ? numero[05][10] - 59 : 59 - numero[05][10];
		diff_pixel[04][06][00] <= numero[06][00] > 121 ? numero[06][00] - 121 : 121 - numero[06][00];
		diff_pixel[04][06][01] <= numero[06][01] > 137 ? numero[06][01] - 137 : 137 - numero[06][01];
		diff_pixel[04][06][02] <= numero[06][02] > 147 ? numero[06][02] - 147 : 147 - numero[06][02];
		diff_pixel[04][06][03] <= numero[06][03] > 140 ? numero[06][03] - 140 : 140 - numero[06][03];
		diff_pixel[04][06][04] <= numero[06][04] > 124 ? numero[06][04] - 124 : 124 - numero[06][04];
		diff_pixel[04][06][05] <= numero[06][05] > 122 ? numero[06][05] - 122 : 122 - numero[06][05];
		diff_pixel[04][06][06] <= numero[06][06] > 140 ? numero[06][06] - 140 : 140 - numero[06][06];
		diff_pixel[04][06][07] <= numero[06][07] > 155 ? numero[06][07] - 155 : 155 - numero[06][07];
		diff_pixel[04][06][08] <= numero[06][08] > 157 ? numero[06][08] - 157 : 157 - numero[06][08];
		diff_pixel[04][06][09] <= numero[06][09] > 130 ? numero[06][09] - 130 : 130 - numero[06][09];
		diff_pixel[04][06][10] <= numero[06][10] > 103 ? numero[06][10] - 103 : 103 - numero[06][10];
		diff_pixel[04][07][00] <= numero[07][00] > 84 ? numero[07][00] - 84 : 84 - numero[07][00];
		diff_pixel[04][07][01] <= numero[07][01] > 103 ? numero[07][01] - 103 : 103 - numero[07][01];
		diff_pixel[04][07][02] <= numero[07][02] > 116 ? numero[07][02] - 116 : 116 - numero[07][02];
		diff_pixel[04][07][03] <= numero[07][03] > 124 ? numero[07][03] - 124 : 124 - numero[07][03];
		diff_pixel[04][07][04] <= numero[07][04] > 124 ? numero[07][04] - 124 : 124 - numero[07][04];
		diff_pixel[04][07][05] <= numero[07][05] > 131 ? numero[07][05] - 131 : 131 - numero[07][05];
		diff_pixel[04][07][06] <= numero[07][06] > 150 ? numero[07][06] - 150 : 150 - numero[07][06];
		diff_pixel[04][07][07] <= numero[07][07] > 161 ? numero[07][07] - 161 : 161 - numero[07][07];
		diff_pixel[04][07][08] <= numero[07][08] > 161 ? numero[07][08] - 161 : 161 - numero[07][08];
		diff_pixel[04][07][09] <= numero[07][09] > 135 ? numero[07][09] - 135 : 135 - numero[07][09];
		diff_pixel[04][07][10] <= numero[07][10] > 106 ? numero[07][10] - 106 : 106 - numero[07][10];
		//diff_pixel[04][08][00] <= numero[08][00] > 0 ? numero[08][00] - 0 : 0 - numero[08][00];
		//diff_pixel[04][08][01] <= numero[08][01] > 0 ? numero[08][01] - 0 : 0 - numero[08][01];
		//diff_pixel[04][08][02] <= numero[08][02] > 0 ? numero[08][02] - 0 : 0 - numero[08][02];
		//diff_pixel[04][08][03] <= numero[08][03] > 0 ? numero[08][03] - 0 : 0 - numero[08][03];
		//diff_pixel[04][08][04] <= numero[08][04] > 4 ? numero[08][04] - 4 : 4 - numero[08][04];
		//diff_pixel[04][08][05] <= numero[08][05] > 33 ? numero[08][05] - 33 : 33 - numero[08][05];
		//diff_pixel[04][08][06] <= numero[08][06] > 83 ? numero[08][06] - 83 : 83 - numero[08][06];
		//diff_pixel[04][08][07] <= numero[08][07] > 118 ? numero[08][07] - 118 : 118 - numero[08][07];
		//diff_pixel[04][08][08] <= numero[08][08] > 122 ? numero[08][08] - 122 : 122 - numero[08][08];
		//diff_pixel[04][08][09] <= numero[08][09] > 91 ? numero[08][09] - 91 : 91 - numero[08][09];
		//diff_pixel[04][08][10] <= numero[08][10] > 43 ? numero[08][10] - 43 : 43 - numero[08][10];
		//diff_pixel[04][09][00] <= numero[09][00] > 0 ? numero[09][00] - 0 : 0 - numero[09][00];
		//diff_pixel[04][09][01] <= numero[09][01] > 0 ? numero[09][01] - 0 : 0 - numero[09][01];
		//diff_pixel[04][09][02] <= numero[09][02] > 0 ? numero[09][02] - 0 : 0 - numero[09][02];
		//diff_pixel[04][09][03] <= numero[09][03] > 0 ? numero[09][03] - 0 : 0 - numero[09][03];
		//diff_pixel[04][09][04] <= numero[09][04] > 3 ? numero[09][04] - 3 : 3 - numero[09][04];
		//diff_pixel[04][09][05] <= numero[09][05] > 31 ? numero[09][05] - 31 : 31 - numero[09][05];
		//diff_pixel[04][09][06] <= numero[09][06] > 83 ? numero[09][06] - 83 : 83 - numero[09][06];
		//diff_pixel[04][09][07] <= numero[09][07] > 119 ? numero[09][07] - 119 : 119 - numero[09][07];
		//diff_pixel[04][09][08] <= numero[09][08] > 126 ? numero[09][08] - 126 : 126 - numero[09][08];
		//diff_pixel[04][09][09] <= numero[09][09] > 97 ? numero[09][09] - 97 : 97 - numero[09][09];
		//diff_pixel[04][09][10] <= numero[09][10] > 48 ? numero[09][10] - 48 : 48 - numero[09][10];
		//diff_pixel[04][10][00] <= numero[10][00] > 0 ? numero[10][00] - 0 : 0 - numero[10][00];
		//diff_pixel[04][10][01] <= numero[10][01] > 0 ? numero[10][01] - 0 : 0 - numero[10][01];
		//diff_pixel[04][10][02] <= numero[10][02] > 0 ? numero[10][02] - 0 : 0 - numero[10][02];
		//diff_pixel[04][10][03] <= numero[10][03] > 0 ? numero[10][03] - 0 : 0 - numero[10][03];
		//diff_pixel[04][10][04] <= numero[10][04] > 4 ? numero[10][04] - 4 : 4 - numero[10][04];
		//diff_pixel[04][10][05] <= numero[10][05] > 24 ? numero[10][05] - 24 : 24 - numero[10][05];
		//diff_pixel[04][10][06] <= numero[10][06] > 58 ? numero[10][06] - 58 : 58 - numero[10][06];
		//diff_pixel[04][10][07] <= numero[10][07] > 82 ? numero[10][07] - 82 : 82 - numero[10][07];
		//diff_pixel[04][10][08] <= numero[10][08] > 83 ? numero[10][08] - 83 : 83 - numero[10][08];
		//diff_pixel[04][10][09] <= numero[10][09] > 62 ? numero[10][09] - 62 : 62 - numero[10][09];
		//diff_pixel[04][10][10] <= numero[10][10] > 29 ? numero[10][10] - 29 : 29 - numero[10][10];
		
		//diff_pixel[05][00][00] <= numero[00][00] > 54 ? numero[00][00] - 54 : 54 - numero[00][00];
		//diff_pixel[05][00][01] <= numero[00][01] > 80 ? numero[00][01] - 80 : 80 - numero[00][01];
		//diff_pixel[05][00][02] <= numero[00][02] > 96 ? numero[00][02] - 96 : 96 - numero[00][02];
		//diff_pixel[05][00][03] <= numero[00][03] > 101 ? numero[00][03] - 101 : 101 - numero[00][03];
		//diff_pixel[05][00][04] <= numero[00][04] > 98 ? numero[00][04] - 98 : 98 - numero[00][04];
		//diff_pixel[05][00][05] <= numero[00][05] > 97 ? numero[00][05] - 97 : 97 - numero[00][05];
		//diff_pixel[05][00][06] <= numero[00][06] > 98 ? numero[00][06] - 98 : 98 - numero[00][06];
		//diff_pixel[05][00][07] <= numero[00][07] > 91 ? numero[00][07] - 91 : 91 - numero[00][07];
		//diff_pixel[05][00][08] <= numero[00][08] > 76 ? numero[00][08] - 76 : 76 - numero[00][08];
		//diff_pixel[05][00][09] <= numero[00][09] > 51 ? numero[00][09] - 51 : 51 - numero[00][09];
		//diff_pixel[05][00][10] <= numero[00][10] > 22 ? numero[00][10] - 22 : 22 - numero[00][10];
		//diff_pixel[05][01][00] <= numero[01][00] > 106 ? numero[01][00] - 106 : 106 - numero[01][00];
		//diff_pixel[05][01][01] <= numero[01][01] > 145 ? numero[01][01] - 145 : 145 - numero[01][01];
		//diff_pixel[05][01][02] <= numero[01][02] > 164 ? numero[01][02] - 164 : 164 - numero[01][02];
		//diff_pixel[05][01][03] <= numero[01][03] > 158 ? numero[01][03] - 158 : 158 - numero[01][03];
		//diff_pixel[05][01][04] <= numero[01][04] > 143 ? numero[01][04] - 143 : 143 - numero[01][04];
		//diff_pixel[05][01][05] <= numero[01][05] > 135 ? numero[01][05] - 135 : 135 - numero[01][05];
		//diff_pixel[05][01][06] <= numero[01][06] > 133 ? numero[01][06] - 133 : 133 - numero[01][06];
		//diff_pixel[05][01][07] <= numero[01][07] > 123 ? numero[01][07] - 123 : 123 - numero[01][07];
		//diff_pixel[05][01][08] <= numero[01][08] > 104 ? numero[01][08] - 104 : 104 - numero[01][08];
		//diff_pixel[05][01][09] <= numero[01][09] > 69 ? numero[01][09] - 69 : 69 - numero[01][09];
		//diff_pixel[05][01][10] <= numero[01][10] > 31 ? numero[01][10] - 31 : 31 - numero[01][10];
		diff_pixel[05][02][00] <= numero[02][00] > 106 ? numero[02][00] - 106 : 106 - numero[02][00];
		diff_pixel[05][02][01] <= numero[02][01] > 133 ? numero[02][01] - 133 : 133 - numero[02][01];
		diff_pixel[05][02][02] <= numero[02][02] > 127 ? numero[02][02] - 127 : 127 - numero[02][02];
		diff_pixel[05][02][03] <= numero[02][03] > 86 ? numero[02][03] - 86 : 86 - numero[02][03];
		diff_pixel[05][02][04] <= numero[02][04] > 41 ? numero[02][04] - 41 : 41 - numero[02][04];
		diff_pixel[05][02][05] <= numero[02][05] > 14 ? numero[02][05] - 14 : 14 - numero[02][05];
		diff_pixel[05][02][06] <= numero[02][06] > 2 ? numero[02][06] - 2 : 2 - numero[02][06];
		diff_pixel[05][02][07] <= numero[02][07] > 2 ? numero[02][07] - 2 : 2 - numero[02][07];
		diff_pixel[05][02][08] <= numero[02][08] > 0 ? numero[02][08] - 0 : 0 - numero[02][08];
		diff_pixel[05][02][09] <= numero[02][09] > 0 ? numero[02][09] - 0 : 0 - numero[02][09];
		diff_pixel[05][02][10] <= numero[02][10] > 0 ? numero[02][10] - 0 : 0 - numero[02][10];
		diff_pixel[05][03][00] <= numero[03][00] > 104 ? numero[03][00] - 104 : 104 - numero[03][00];
		diff_pixel[05][03][01] <= numero[03][01] > 143 ? numero[03][01] - 143 : 143 - numero[03][01];
		diff_pixel[05][03][02] <= numero[03][02] > 155 ? numero[03][02] - 155 : 155 - numero[03][02];
		diff_pixel[05][03][03] <= numero[03][03] > 144 ? numero[03][03] - 144 : 144 - numero[03][03];
		diff_pixel[05][03][04] <= numero[03][04] > 125 ? numero[03][04] - 125 : 125 - numero[03][04];
		diff_pixel[05][03][05] <= numero[03][05] > 113 ? numero[03][05] - 113 : 113 - numero[03][05];
		diff_pixel[05][03][06] <= numero[03][06] > 112 ? numero[03][06] - 112 : 112 - numero[03][06];
		diff_pixel[05][03][07] <= numero[03][07] > 105 ? numero[03][07] - 105 : 105 - numero[03][07];
		diff_pixel[05][03][08] <= numero[03][08] > 89 ? numero[03][08] - 89 : 89 - numero[03][08];
		diff_pixel[05][03][09] <= numero[03][09] > 60 ? numero[03][09] - 60 : 60 - numero[03][09];
		diff_pixel[05][03][10] <= numero[03][10] > 33 ? numero[03][10] - 33 : 33 - numero[03][10];
		diff_pixel[05][04][00] <= numero[04][00] > 73 ? numero[04][00] - 73 : 73 - numero[04][00];
		diff_pixel[05][04][01] <= numero[04][01] > 107 ? numero[04][01] - 107 : 107 - numero[04][01];
		diff_pixel[05][04][02] <= numero[04][02] > 122 ? numero[04][02] - 122 : 122 - numero[04][02];
		diff_pixel[05][04][03] <= numero[04][03] > 128 ? numero[04][03] - 128 : 128 - numero[04][03];
		diff_pixel[05][04][04] <= numero[04][04] > 122 ? numero[04][04] - 122 : 122 - numero[04][04];
		diff_pixel[05][04][05] <= numero[04][05] > 123 ? numero[04][05] - 123 : 123 - numero[04][05];
		diff_pixel[05][04][06] <= numero[04][06] > 128 ? numero[04][06] - 128 : 128 - numero[04][06];
		diff_pixel[05][04][07] <= numero[04][07] > 132 ? numero[04][07] - 132 : 132 - numero[04][07];
		diff_pixel[05][04][08] <= numero[04][08] > 123 ? numero[04][08] - 123 : 123 - numero[04][08];
		diff_pixel[05][04][09] <= numero[04][09] > 98 ? numero[04][09] - 98 : 98 - numero[04][09];
		diff_pixel[05][04][10] <= numero[04][10] > 69 ? numero[04][10] - 69 : 69 - numero[04][10];
		diff_pixel[05][05][00] <= numero[05][00] > 0 ? numero[05][00] - 0 : 0 - numero[05][00];
		diff_pixel[05][05][01] <= numero[05][01] > 7 ? numero[05][01] - 7 : 7 - numero[05][01];
		diff_pixel[05][05][02] <= numero[05][02] > 5 ? numero[05][02] - 5 : 5 - numero[05][02];
		diff_pixel[05][05][03] <= numero[05][03] > 6 ? numero[05][03] - 6 : 6 - numero[05][03];
		diff_pixel[05][05][04] <= numero[05][04] > 2 ? numero[05][04] - 2 : 2 - numero[05][04];
		diff_pixel[05][05][05] <= numero[05][05] > 8 ? numero[05][05] - 8 : 8 - numero[05][05];
		diff_pixel[05][05][06] <= numero[05][06] > 29 ? numero[05][06] - 29 : 29 - numero[05][06];
		diff_pixel[05][05][07] <= numero[05][07] > 64 ? numero[05][07] - 64 : 64 - numero[05][07];
		diff_pixel[05][05][08] <= numero[05][08] > 106 ? numero[05][08] - 106 : 106 - numero[05][08];
		diff_pixel[05][05][09] <= numero[05][09] > 118 ? numero[05][09] - 118 : 118 - numero[05][09];
		diff_pixel[05][05][10] <= numero[05][10] > 120 ? numero[05][10] - 120 : 120 - numero[05][10];
		diff_pixel[05][06][00] <= numero[06][00] > 1 ? numero[06][00] - 1 : 1 - numero[06][00];
		diff_pixel[05][06][01] <= numero[06][01] > 0 ? numero[06][01] - 0 : 0 - numero[06][01];
		diff_pixel[05][06][02] <= numero[06][02] > 0 ? numero[06][02] - 0 : 0 - numero[06][02];
		diff_pixel[05][06][03] <= numero[06][03] > 0 ? numero[06][03] - 0 : 0 - numero[06][03];
		diff_pixel[05][06][04] <= numero[06][04] > 0 ? numero[06][04] - 0 : 0 - numero[06][04];
		diff_pixel[05][06][05] <= numero[06][05] > 0 ? numero[06][05] - 0 : 0 - numero[06][05];
		diff_pixel[05][06][06] <= numero[06][06] > 24 ? numero[06][06] - 24 : 24 - numero[06][06];
		diff_pixel[05][06][07] <= numero[06][07] > 61 ? numero[06][07] - 61 : 61 - numero[06][07];
		diff_pixel[05][06][08] <= numero[06][08] > 109 ? numero[06][08] - 109 : 109 - numero[06][08];
		diff_pixel[05][06][09] <= numero[06][09] > 126 ? numero[06][09] - 126 : 126 - numero[06][09];
		diff_pixel[05][06][10] <= numero[06][10] > 125 ? numero[06][10] - 125 : 125 - numero[06][10];
		diff_pixel[05][07][00] <= numero[07][00] > 42 ? numero[07][00] - 42 : 42 - numero[07][00];
		diff_pixel[05][07][01] <= numero[07][01] > 37 ? numero[07][01] - 37 : 37 - numero[07][01];
		diff_pixel[05][07][02] <= numero[07][02] > 31 ? numero[07][02] - 31 : 31 - numero[07][02];
		diff_pixel[05][07][03] <= numero[07][03] > 19 ? numero[07][03] - 19 : 19 - numero[07][03];
		diff_pixel[05][07][04] <= numero[07][04] > 3 ? numero[07][04] - 3 : 3 - numero[07][04];
		diff_pixel[05][07][05] <= numero[07][05] > 0 ? numero[07][05] - 0 : 0 - numero[07][05];
		diff_pixel[05][07][06] <= numero[07][06] > 22 ? numero[07][06] - 22 : 22 - numero[07][06];
		diff_pixel[05][07][07] <= numero[07][07] > 59 ? numero[07][07] - 59 : 59 - numero[07][07];
		diff_pixel[05][07][08] <= numero[07][08] > 106 ? numero[07][08] - 106 : 106 - numero[07][08];
		diff_pixel[05][07][09] <= numero[07][09] > 122 ? numero[07][09] - 122 : 122 - numero[07][09];
		diff_pixel[05][07][10] <= numero[07][10] > 120 ? numero[07][10] - 120 : 120 - numero[07][10];
		//diff_pixel[05][08][00] <= numero[08][00] > 99 ? numero[08][00] - 99 : 99 - numero[08][00];
		//diff_pixel[05][08][01] <= numero[08][01] > 125 ? numero[08][01] - 125 : 125 - numero[08][01];
		//diff_pixel[05][08][02] <= numero[08][02] > 120 ? numero[08][02] - 120 : 120 - numero[08][02];
		//diff_pixel[05][08][03] <= numero[08][03] > 78 ? numero[08][03] - 78 : 78 - numero[08][03];
		//diff_pixel[05][08][04] <= numero[08][04] > 28 ? numero[08][04] - 28 : 28 - numero[08][04];
		//diff_pixel[05][08][05] <= numero[08][05] > 4 ? numero[08][05] - 4 : 4 - numero[08][05];
		//diff_pixel[05][08][06] <= numero[08][06] > 21 ? numero[08][06] - 21 : 21 - numero[08][06];
		//diff_pixel[05][08][07] <= numero[08][07] > 61 ? numero[08][07] - 61 : 61 - numero[08][07];
		//diff_pixel[05][08][08] <= numero[08][08] > 116 ? numero[08][08] - 116 : 116 - numero[08][08];
		//diff_pixel[05][08][09] <= numero[08][09] > 133 ? numero[08][09] - 133 : 133 - numero[08][09];
		//diff_pixel[05][08][10] <= numero[08][10] > 121 ? numero[08][10] - 121 : 121 - numero[08][10];
		//diff_pixel[05][09][00] <= numero[09][00] > 52 ? numero[09][00] - 52 : 52 - numero[09][00];
		//diff_pixel[05][09][01] <= numero[09][01] > 92 ? numero[09][01] - 92 : 92 - numero[09][01];
		//diff_pixel[05][09][02] <= numero[09][02] > 131 ? numero[09][02] - 131 : 131 - numero[09][02];
		//diff_pixel[05][09][03] <= numero[09][03] > 139 ? numero[09][03] - 139 : 139 - numero[09][03];
		//diff_pixel[05][09][04] <= numero[09][04] > 137 ? numero[09][04] - 137 : 137 - numero[09][04];
		//diff_pixel[05][09][05] <= numero[09][05] > 132 ? numero[09][05] - 132 : 132 - numero[09][05];
		//diff_pixel[05][09][06] <= numero[09][06] > 134 ? numero[09][06] - 134 : 134 - numero[09][06];
		//diff_pixel[05][09][07] <= numero[09][07] > 136 ? numero[09][07] - 136 : 136 - numero[09][07];
		//diff_pixel[05][09][08] <= numero[09][08] > 134 ? numero[09][08] - 134 : 134 - numero[09][08];
		//diff_pixel[05][09][09] <= numero[09][09] > 109 ? numero[09][09] - 109 : 109 - numero[09][09];
		//diff_pixel[05][09][10] <= numero[09][10] > 67 ? numero[09][10] - 67 : 67 - numero[09][10];
		//diff_pixel[05][10][00] <= numero[10][00] > 15 ? numero[10][00] - 15 : 15 - numero[10][00];
		//diff_pixel[05][10][01] <= numero[10][01] > 47 ? numero[10][01] - 47 : 47 - numero[10][01];
		//diff_pixel[05][10][02] <= numero[10][02] > 82 ? numero[10][02] - 82 : 82 - numero[10][02];
		//diff_pixel[05][10][03] <= numero[10][03] > 105 ? numero[10][03] - 105 : 105 - numero[10][03];
		//diff_pixel[05][10][04] <= numero[10][04] > 115 ? numero[10][04] - 115 : 115 - numero[10][04];
		//diff_pixel[05][10][05] <= numero[10][05] > 116 ? numero[10][05] - 116 : 116 - numero[10][05];
		//diff_pixel[05][10][06] <= numero[10][06] > 119 ? numero[10][06] - 119 : 119 - numero[10][06];
		//diff_pixel[05][10][07] <= numero[10][07] > 108 ? numero[10][07] - 108 : 108 - numero[10][07];
		//diff_pixel[05][10][08] <= numero[10][08] > 95 ? numero[10][08] - 95 : 95 - numero[10][08];
		//diff_pixel[05][10][09] <= numero[10][09] > 64 ? numero[10][09] - 64 : 64 - numero[10][09];
//		
		//diff_pixel[06][00][00] <= numero[00][00] > 19 ? numero[00][00] - 19 : 19 - numero[00][00];
		//diff_pixel[06][00][01] <= numero[00][01] > 30 ? numero[00][01] - 30 : 30 - numero[00][01];
		//diff_pixel[06][00][02] <= numero[00][02] > 41 ? numero[00][02] - 41 : 41 - numero[00][02];
		//diff_pixel[06][00][03] <= numero[00][03] > 69 ? numero[00][03] - 69 : 69 - numero[00][03];
		//diff_pixel[06][00][04] <= numero[00][04] > 84 ? numero[00][04] - 84 : 84 - numero[00][04];
		//diff_pixel[06][00][05] <= numero[00][05] > 100 ? numero[00][05] - 100 : 100 - numero[00][05];
		//diff_pixel[06][00][06] <= numero[00][06] > 104 ? numero[00][06] - 104 : 104 - numero[00][06];
		//diff_pixel[06][00][07] <= numero[00][07] > 96 ? numero[00][07] - 96 : 96 - numero[00][07];
		//diff_pixel[06][00][08] <= numero[00][08] > 73 ? numero[00][08] - 73 : 73 - numero[00][08];
		//diff_pixel[06][00][09] <= numero[00][09] > 48 ? numero[00][09] - 48 : 48 - numero[00][09];
		//diff_pixel[06][00][10] <= numero[00][10] > 21 ? numero[00][10] - 21 : 21 - numero[00][10];
		//diff_pixel[06][01][00] <= numero[01][00] > 9 ? numero[01][00] - 9 : 9 - numero[01][00];
		//diff_pixel[06][01][01] <= numero[01][01] > 35 ? numero[01][01] - 35 : 35 - numero[01][01];
		//diff_pixel[06][01][02] <= numero[01][02] > 70 ? numero[01][02] - 70 : 70 - numero[01][02];
		//diff_pixel[06][01][03] <= numero[01][03] > 111 ? numero[01][03] - 111 : 111 - numero[01][03];
		//diff_pixel[06][01][04] <= numero[01][04] > 136 ? numero[01][04] - 136 : 136 - numero[01][04];
		//diff_pixel[06][01][05] <= numero[01][05] > 143 ? numero[01][05] - 143 : 143 - numero[01][05];
		//diff_pixel[06][01][06] <= numero[01][06] > 142 ? numero[01][06] - 142 : 142 - numero[01][06];
		//diff_pixel[06][01][07] <= numero[01][07] > 125 ? numero[01][07] - 125 : 125 - numero[01][07];
		//diff_pixel[06][01][08] <= numero[01][08] > 102 ? numero[01][08] - 102 : 102 - numero[01][08];
		//diff_pixel[06][01][09] <= numero[01][09] > 70 ? numero[01][09] - 70 : 70 - numero[01][09];
		//diff_pixel[06][01][10] <= numero[01][10] > 32 ? numero[01][10] - 32 : 32 - numero[01][10];
		diff_pixel[06][02][00] <= numero[02][00] > 44 ? numero[02][00] - 44 : 44 - numero[02][00];
		diff_pixel[06][02][01] <= numero[02][01] > 72 ? numero[02][01] - 72 : 72 - numero[02][01];
		diff_pixel[06][02][02] <= numero[02][02] > 111 ? numero[02][02] - 111 : 111 - numero[02][02];
		diff_pixel[06][02][03] <= numero[02][03] > 126 ? numero[02][03] - 126 : 126 - numero[02][03];
		diff_pixel[06][02][04] <= numero[02][04] > 106 ? numero[02][04] - 106 : 106 - numero[02][04];
		diff_pixel[06][02][05] <= numero[02][05] > 59 ? numero[02][05] - 59 : 59 - numero[02][05];
		diff_pixel[06][02][06] <= numero[02][06] > 23 ? numero[02][06] - 23 : 23 - numero[02][06];
		diff_pixel[06][02][07] <= numero[02][07] > 2 ? numero[02][07] - 2 : 2 - numero[02][07];
		diff_pixel[06][02][08] <= numero[02][08] > 0 ? numero[02][08] - 0 : 0 - numero[02][08];
		diff_pixel[06][02][09] <= numero[02][09] > 0 ? numero[02][09] - 0 : 0 - numero[02][09];
		diff_pixel[06][02][10] <= numero[02][10] > 0 ? numero[02][10] - 0 : 0 - numero[02][10];
		diff_pixel[06][03][00] <= numero[03][00] > 100 ? numero[03][00] - 100 : 100 - numero[03][00];
		diff_pixel[06][03][01] <= numero[03][01] > 111 ? numero[03][01] - 111 : 111 - numero[03][01];
		diff_pixel[06][03][02] <= numero[03][02] > 120 ? numero[03][02] - 120 : 120 - numero[03][02];
		diff_pixel[06][03][03] <= numero[03][03] > 100 ? numero[03][03] - 100 : 100 - numero[03][03];
		diff_pixel[06][03][04] <= numero[03][04] > 59 ? numero[03][04] - 59 : 59 - numero[03][04];
		diff_pixel[06][03][05] <= numero[03][05] > 21 ? numero[03][05] - 21 : 21 - numero[03][05];
		diff_pixel[06][03][06] <= numero[03][06] > 0 ? numero[03][06] - 0 : 0 - numero[03][06];
		diff_pixel[06][03][07] <= numero[03][07] > 0 ? numero[03][07] - 0 : 0 - numero[03][07];
		diff_pixel[06][03][08] <= numero[03][08] > 0 ? numero[03][08] - 0 : 0 - numero[03][08];
		diff_pixel[06][03][09] <= numero[03][09] > 0 ? numero[03][09] - 0 : 0 - numero[03][09];
		diff_pixel[06][03][10] <= numero[03][10] > 0 ? numero[03][10] - 0 : 0 - numero[03][10];
		diff_pixel[06][04][00] <= numero[04][00] > 119 ? numero[04][00] - 119 : 119 - numero[04][00];
		diff_pixel[06][04][01] <= numero[04][01] > 129 ? numero[04][01] - 129 : 129 - numero[04][01];
		diff_pixel[06][04][02] <= numero[04][02] > 129 ? numero[04][02] - 129 : 129 - numero[04][02];
		diff_pixel[06][04][03] <= numero[04][03] > 107 ? numero[04][03] - 107 : 107 - numero[04][03];
		diff_pixel[06][04][04] <= numero[04][04] > 73 ? numero[04][04] - 73 : 73 - numero[04][04];
		diff_pixel[06][04][05] <= numero[04][05] > 53 ? numero[04][05] - 53 : 53 - numero[04][05];
		diff_pixel[06][04][06] <= numero[04][06] > 45 ? numero[04][06] - 45 : 45 - numero[04][06];
		diff_pixel[06][04][07] <= numero[04][07] > 43 ? numero[04][07] - 43 : 43 - numero[04][07];
		diff_pixel[06][04][08] <= numero[04][08] > 36 ? numero[04][08] - 36 : 36 - numero[04][08];
		diff_pixel[06][04][09] <= numero[04][09] > 21 ? numero[04][09] - 21 : 21 - numero[04][09];
		diff_pixel[06][04][10] <= numero[04][10] > 15 ? numero[04][10] - 15 : 15 - numero[04][10];
		diff_pixel[06][05][00] <= numero[05][00] > 126 ? numero[05][00] - 126 : 126 - numero[05][00];
		diff_pixel[06][05][01] <= numero[05][01] > 148 ? numero[05][01] - 148 : 148 - numero[05][01];
		diff_pixel[06][05][02] <= numero[05][02] > 170 ? numero[05][02] - 170 : 170 - numero[05][02];
		diff_pixel[06][05][03] <= numero[05][03] > 179 ? numero[05][03] - 179 : 179 - numero[05][03];
		diff_pixel[06][05][04] <= numero[05][04] > 174 ? numero[05][04] - 174 : 174 - numero[05][04];
		diff_pixel[06][05][05] <= numero[05][05] > 168 ? numero[05][05] - 168 : 168 - numero[05][05];
		diff_pixel[06][05][06] <= numero[05][06] > 168 ? numero[05][06] - 168 : 168 - numero[05][06];
		diff_pixel[06][05][07] <= numero[05][07] > 157 ? numero[05][07] - 157 : 157 - numero[05][07];
		diff_pixel[06][05][08] <= numero[05][08] > 129 ? numero[05][08] - 129 : 129 - numero[05][08];
		diff_pixel[06][05][09] <= numero[05][09] > 86 ? numero[05][09] - 86 : 86 - numero[05][09];
		diff_pixel[06][05][10] <= numero[05][10] > 48 ? numero[05][10] - 48 : 48 - numero[05][10];
		diff_pixel[06][06][00] <= numero[06][00] > 122 ? numero[06][00] - 122 : 122 - numero[06][00];
		diff_pixel[06][06][01] <= numero[06][01] > 134 ? numero[06][01] - 134 : 134 - numero[06][01];
		diff_pixel[06][06][02] <= numero[06][02] > 136 ? numero[06][02] - 136 : 136 - numero[06][02];
		diff_pixel[06][06][03] <= numero[06][03] > 117 ? numero[06][03] - 117 : 117 - numero[06][03];
		diff_pixel[06][06][04] <= numero[06][04] > 86 ? numero[06][04] - 86 : 86 - numero[06][04];
		diff_pixel[06][06][05] <= numero[06][05] > 71 ? numero[06][05] - 71 : 71 - numero[06][05];
		diff_pixel[06][06][06] <= numero[06][06] > 81 ? numero[06][06] - 81 : 81 - numero[06][06];
		diff_pixel[06][06][07] <= numero[06][07] > 101 ? numero[06][07] - 101 : 101 - numero[06][07];
		diff_pixel[06][06][08] <= numero[06][08] > 124 ? numero[06][08] - 124 : 124 - numero[06][08];
		diff_pixel[06][06][09] <= numero[06][09] > 117 ? numero[06][09] - 117 : 117 - numero[06][09];
		diff_pixel[06][06][10] <= numero[06][10] > 99 ? numero[06][10] - 99 : 99 - numero[06][10];
		diff_pixel[06][07][00] <= numero[07][00] > 115 ? numero[07][00] - 115 : 115 - numero[07][00];
		diff_pixel[06][07][01] <= numero[07][01] > 126 ? numero[07][01] - 126 : 126 - numero[07][01];
		diff_pixel[06][07][02] <= numero[07][02] > 118 ? numero[07][02] - 118 : 118 - numero[07][02];
		diff_pixel[06][07][03] <= numero[07][03] > 80 ? numero[07][03] - 80 : 80 - numero[07][03];
		diff_pixel[06][07][04] <= numero[07][04] > 33 ? numero[07][04] - 33 : 33 - numero[07][04];
		diff_pixel[06][07][05] <= numero[07][05] > 9 ? numero[07][05] - 9 : 9 - numero[07][05];
		diff_pixel[06][07][06] <= numero[07][06] > 20 ? numero[07][06] - 20 : 20 - numero[07][06];
		diff_pixel[06][07][07] <= numero[07][07] > 60 ? numero[07][07] - 60 : 60 - numero[07][07];
		diff_pixel[06][07][08] <= numero[07][08] > 108 ? numero[07][08] - 108 : 108 - numero[07][08];
		diff_pixel[06][07][09] <= numero[07][09] > 125 ? numero[07][09] - 125 : 125 - numero[07][09];
		diff_pixel[06][07][10] <= numero[07][10] > 119 ? numero[07][10] - 119 : 119 - numero[07][10];
		//diff_pixel[06][08][00] <= numero[08][00] > 105 ? numero[08][00] - 105 : 105 - numero[08][00];
		//diff_pixel[06][08][01] <= numero[08][01] > 131 ? numero[08][01] - 131 : 131 - numero[08][01];
		//diff_pixel[06][08][02] <= numero[08][02] > 120 ? numero[08][02] - 120 : 120 - numero[08][02];
		//diff_pixel[06][08][03] <= numero[08][03] > 78 ? numero[08][03] - 78 : 78 - numero[08][03];
		//diff_pixel[06][08][04] <= numero[08][04] > 28 ? numero[08][04] - 28 : 28 - numero[08][04];
		//diff_pixel[06][08][05] <= numero[08][05] > 4 ? numero[08][05] - 4 : 4 - numero[08][05];
		//diff_pixel[06][08][06] <= numero[08][06] > 22 ? numero[08][06] - 22 : 22 - numero[08][06];
		//diff_pixel[06][08][07] <= numero[08][07] > 62 ? numero[08][07] - 62 : 62 - numero[08][07];
		//diff_pixel[06][08][08] <= numero[08][08] > 115 ? numero[08][08] - 115 : 115 - numero[08][08];
		//diff_pixel[06][08][09] <= numero[08][09] > 134 ? numero[08][09] - 134 : 134 - numero[08][09];
		//diff_pixel[06][08][10] <= numero[08][10] > 118 ? numero[08][10] - 118 : 118 - numero[08][10];
		//diff_pixel[06][09][00] <= numero[09][00] > 58 ? numero[09][00] - 58 : 58 - numero[09][00];
		//diff_pixel[06][09][01] <= numero[09][01] > 95 ? numero[09][01] - 95 : 95 - numero[09][01];
		//diff_pixel[06][09][02] <= numero[09][02] > 131 ? numero[09][02] - 131 : 131 - numero[09][02];
		//diff_pixel[06][09][03] <= numero[09][03] > 142 ? numero[09][03] - 142 : 142 - numero[09][03];
		//diff_pixel[06][09][04] <= numero[09][04] > 138 ? numero[09][04] - 138 : 138 - numero[09][04];
		//diff_pixel[06][09][05] <= numero[09][05] > 134 ? numero[09][05] - 134 : 134 - numero[09][05];
		//diff_pixel[06][09][06] <= numero[09][06] > 134 ? numero[09][06] - 134 : 134 - numero[09][06];
		//diff_pixel[06][09][07] <= numero[09][07] > 136 ? numero[09][07] - 136 : 136 - numero[09][07];
		//diff_pixel[06][09][08] <= numero[09][08] > 134 ? numero[09][08] - 134 : 134 - numero[09][08];
		//diff_pixel[06][09][09] <= numero[09][09] > 110 ? numero[09][09] - 110 : 110 - numero[09][09];
		//diff_pixel[06][09][10] <= numero[09][10] > 66 ? numero[09][10] - 66 : 66 - numero[09][10];
		//diff_pixel[06][10][00] <= numero[10][00] > 16 ? numero[10][00] - 16 : 16 - numero[10][00];
		//diff_pixel[06][10][01] <= numero[10][01] > 47 ? numero[10][01] - 47 : 47 - numero[10][01];
		//diff_pixel[06][10][02] <= numero[10][02] > 80 ? numero[10][02] - 80 : 80 - numero[10][02];
		//diff_pixel[06][10][03] <= numero[10][03] > 103 ? numero[10][03] - 103 : 103 - numero[10][03];
		//diff_pixel[06][10][04] <= numero[10][04] > 113 ? numero[10][04] - 113 : 113 - numero[10][04];
		//diff_pixel[06][10][05] <= numero[10][05] > 115 ? numero[10][05] - 115 : 115 - numero[10][05];
		//diff_pixel[06][10][06] <= numero[10][06] > 119 ? numero[10][06] - 119 : 119 - numero[10][06];
		//diff_pixel[06][10][07] <= numero[10][07] > 108 ? numero[10][07] - 108 : 108 - numero[10][07];
		//diff_pixel[06][10][08] <= numero[10][08] > 95 ? numero[10][08] - 95 : 95 - numero[10][08];
		//diff_pixel[06][10][09] <= numero[10][09] > 64 ? numero[10][09] - 64 : 64 - numero[10][09];
		//diff_pixel[06][10][10] <= numero[10][10] > 30 ? numero[10][10] - 30 : 30 - numero[10][10];
		
		//diff_pixel[07][00][00] <= numero[00][00] > 54 ? numero[00][00] - 54 : 54 - numero[00][00];
		//diff_pixel[07][00][01] <= numero[00][01] > 80 ? numero[00][01] - 80 : 80 - numero[00][01];
		//diff_pixel[07][00][02] <= numero[00][02] > 95 ? numero[00][02] - 95 : 95 - numero[00][02];
		//diff_pixel[07][00][03] <= numero[00][03] > 100 ? numero[00][03] - 100 : 100 - numero[00][03];
		//diff_pixel[07][00][04] <= numero[00][04] > 95 ? numero[00][04] - 95 : 95 - numero[00][04];
		//diff_pixel[07][00][05] <= numero[00][05] > 94 ? numero[00][05] - 94 : 94 - numero[00][05];
		//diff_pixel[07][00][06] <= numero[00][06] > 97 ? numero[00][06] - 97 : 97 - numero[00][06];
		//diff_pixel[07][00][07] <= numero[00][07] > 97 ? numero[00][07] - 97 : 97 - numero[00][07];
		//diff_pixel[07][00][08] <= numero[00][08] > 96 ? numero[00][08] - 96 : 96 - numero[00][08];
		//diff_pixel[07][00][09] <= numero[00][09] > 83 ? numero[00][09] - 83 : 83 - numero[00][09];
		//diff_pixel[07][00][10] <= numero[00][10] > 66 ? numero[00][10] - 66 : 66 - numero[00][10];
		//diff_pixel[07][01][00] <= numero[01][00] > 104 ? numero[01][00] - 104 : 104 - numero[01][00];
		//diff_pixel[07][01][01] <= numero[01][01] > 146 ? numero[01][01] - 146 : 146 - numero[01][01];
		//diff_pixel[07][01][02] <= numero[01][02] > 161 ? numero[01][02] - 161 : 161 - numero[01][02];
		//diff_pixel[07][01][03] <= numero[01][03] > 156 ? numero[01][03] - 156 : 156 - numero[01][03];
		//diff_pixel[07][01][04] <= numero[01][04] > 139 ? numero[01][04] - 139 : 139 - numero[01][04];
		//diff_pixel[07][01][05] <= numero[01][05] > 132 ? numero[01][05] - 132 : 132 - numero[01][05];
		//diff_pixel[07][01][06] <= numero[01][06] > 136 ? numero[01][06] - 136 : 136 - numero[01][06];
		//diff_pixel[07][01][07] <= numero[01][07] > 147 ? numero[01][07] - 147 : 147 - numero[01][07];
		//diff_pixel[07][01][08] <= numero[01][08] > 159 ? numero[01][08] - 159 : 159 - numero[01][08];
		//diff_pixel[07][01][09] <= numero[01][09] > 146 ? numero[01][09] - 146 : 146 - numero[01][09];
		//diff_pixel[07][01][10] <= numero[01][10] > 120 ? numero[01][10] - 120 : 120 - numero[01][10];
		diff_pixel[07][02][00] <= numero[02][00] > 108 ? numero[02][00] - 108 : 108 - numero[02][00];
		diff_pixel[07][02][01] <= numero[02][01] > 131 ? numero[02][01] - 131 : 131 - numero[02][01];
		diff_pixel[07][02][02] <= numero[02][02] > 126 ? numero[02][02] - 126 : 126 - numero[02][02];
		diff_pixel[07][02][03] <= numero[02][03] > 87 ? numero[02][03] - 87 : 87 - numero[02][03];
		diff_pixel[07][02][04] <= numero[02][04] > 38 ? numero[02][04] - 38 : 38 - numero[02][04];
		diff_pixel[07][02][05] <= numero[02][05] > 16 ? numero[02][05] - 16 : 16 - numero[02][05];
		diff_pixel[07][02][06] <= numero[02][06] > 28 ? numero[02][06] - 28 : 28 - numero[02][06];
		diff_pixel[07][02][07] <= numero[02][07] > 66 ? numero[02][07] - 66 : 66 - numero[02][07];
		diff_pixel[07][02][08] <= numero[02][08] > 115 ? numero[02][08] - 115 : 115 - numero[02][08];
		diff_pixel[07][02][09] <= numero[02][09] > 131 ? numero[02][09] - 131 : 131 - numero[02][09];
		diff_pixel[07][02][10] <= numero[02][10] > 115 ? numero[02][10] - 115 : 115 - numero[02][10];
		diff_pixel[07][03][00] <= numero[03][00] > 31 ? numero[03][00] - 31 : 31 - numero[03][00];
		diff_pixel[07][03][01] <= numero[03][01] > 43 ? numero[03][01] - 43 : 43 - numero[03][01];
		diff_pixel[07][03][02] <= numero[03][02] > 38 ? numero[03][02] - 38 : 38 - numero[03][02];
		diff_pixel[07][03][03] <= numero[03][03] > 22 ? numero[03][03] - 22 : 22 - numero[03][03];
		diff_pixel[07][03][04] <= numero[03][04] > 12 ? numero[03][04] - 12 : 12 - numero[03][04];
		diff_pixel[07][03][05] <= numero[03][05] > 21 ? numero[03][05] - 21 : 21 - numero[03][05];
		diff_pixel[07][03][06] <= numero[03][06] > 60 ? numero[03][06] - 60 : 60 - numero[03][06];
		diff_pixel[07][03][07] <= numero[03][07] > 99 ? numero[03][07] - 99 : 99 - numero[03][07];
		diff_pixel[07][03][08] <= numero[03][08] > 123 ? numero[03][08] - 123 : 123 - numero[03][08];
		diff_pixel[07][03][09] <= numero[03][09] > 111 ? numero[03][09] - 111 : 111 - numero[03][09];
		diff_pixel[07][03][10] <= numero[03][10] > 82 ? numero[03][10] - 82 : 82 - numero[03][10];
		diff_pixel[07][04][00] <= numero[04][00] > 0 ? numero[04][00] - 0 : 0 - numero[04][00];
		diff_pixel[07][04][01] <= numero[04][01] > 0 ? numero[04][01] - 0 : 0 - numero[04][01];
		diff_pixel[07][04][02] <= numero[04][02] > 0 ? numero[04][02] - 0 : 0 - numero[04][02];
		diff_pixel[07][04][03] <= numero[04][03] > 5 ? numero[04][03] - 5 : 5 - numero[04][03];
		diff_pixel[07][04][04] <= numero[04][04] > 30 ? numero[04][04] - 30 : 30 - numero[04][04];
		diff_pixel[07][04][05] <= numero[04][05] > 65 ? numero[04][05] - 65 : 65 - numero[04][05];
		diff_pixel[07][04][06] <= numero[04][06] > 101 ? numero[04][06] - 101 : 101 - numero[04][06];
		diff_pixel[07][04][07] <= numero[04][07] > 122 ? numero[04][07] - 122 : 122 - numero[04][07];
		diff_pixel[07][04][08] <= numero[04][08] > 109 ? numero[04][08] - 109 : 109 - numero[04][08];
		diff_pixel[07][04][09] <= numero[04][09] > 72 ? numero[04][09] - 72 : 72 - numero[04][09];
		diff_pixel[07][04][10] <= numero[04][10] > 37 ? numero[04][10] - 37 : 37 - numero[04][10];
		diff_pixel[07][05][00] <= numero[05][00] > 0 ? numero[05][00] - 0 : 0 - numero[05][00];
		diff_pixel[07][05][01] <= numero[05][01] > 0 ? numero[05][01] - 0 : 0 - numero[05][01];
		diff_pixel[07][05][02] <= numero[05][02] > 0 ? numero[05][02] - 0 : 0 - numero[05][02];
		diff_pixel[07][05][03] <= numero[05][03] > 20 ? numero[05][03] - 20 : 20 - numero[05][03];
		diff_pixel[07][05][04] <= numero[05][04] > 62 ? numero[05][04] - 62 : 62 - numero[05][04];
		diff_pixel[07][05][05] <= numero[05][05] > 108 ? numero[05][05] - 108 : 108 - numero[05][05];
		diff_pixel[07][05][06] <= numero[05][06] > 129 ? numero[05][06] - 129 : 129 - numero[05][06];
		diff_pixel[07][05][07] <= numero[05][07] > 115 ? numero[05][07] - 115 : 115 - numero[05][07];
		diff_pixel[07][05][08] <= numero[05][08] > 71 ? numero[05][08] - 71 : 71 - numero[05][08];
		diff_pixel[07][05][09] <= numero[05][09] > 25 ? numero[05][09] - 25 : 25 - numero[05][09];
		diff_pixel[07][05][10] <= numero[05][10] > 7 ? numero[05][10] - 7 : 7 - numero[05][10];
		diff_pixel[07][06][00] <= numero[06][00] > 9 ? numero[06][00] - 9 : 9 - numero[06][00];
		diff_pixel[07][06][01] <= numero[06][01] > 3 ? numero[06][01] - 3 : 3 - numero[06][01];
		diff_pixel[07][06][02] <= numero[06][02] > 28 ? numero[06][02] - 28 : 28 - numero[06][02];
		diff_pixel[07][06][03] <= numero[06][03] > 75 ? numero[06][03] - 75 : 75 - numero[06][03];
		diff_pixel[07][06][04] <= numero[06][04] > 110 ? numero[06][04] - 110 : 110 - numero[06][04];
		diff_pixel[07][06][05] <= numero[06][05] > 126 ? numero[06][05] - 126 : 126 - numero[06][05];
		diff_pixel[07][06][06] <= numero[06][06] > 106 ? numero[06][06] - 106 : 106 - numero[06][06];
		diff_pixel[07][06][07] <= numero[06][07] > 68 ? numero[06][07] - 68 : 68 - numero[06][07];
		diff_pixel[07][06][08] <= numero[06][08] > 27 ? numero[06][08] - 27 : 27 - numero[06][08];
		diff_pixel[07][06][09] <= numero[06][09] > 0 ? numero[06][09] - 0 : 0 - numero[06][09];
		diff_pixel[07][06][10] <= numero[06][10] > 0 ? numero[06][10] - 0 : 0 - numero[06][10];
		diff_pixel[07][07][00] <= numero[07][00] > 3 ? numero[07][00] - 3 : 3 - numero[07][00];
		diff_pixel[07][07][01] <= numero[07][01] > 6 ? numero[07][01] - 6 : 6 - numero[07][01];
		diff_pixel[07][07][02] <= numero[07][02] > 42 ? numero[07][02] - 42 : 42 - numero[07][02];
		diff_pixel[07][07][03] <= numero[07][03] > 98 ? numero[07][03] - 98 : 98 - numero[07][03];
		diff_pixel[07][07][04] <= numero[07][04] > 130 ? numero[07][04] - 130 : 130 - numero[07][04];
		diff_pixel[07][07][05] <= numero[07][05] > 129 ? numero[07][05] - 129 : 129 - numero[07][05];
		diff_pixel[07][07][06] <= numero[07][06] > 91 ? numero[07][06] - 91 : 91 - numero[07][06];
		diff_pixel[07][07][07] <= numero[07][07] > 40 ? numero[07][07] - 40 : 40 - numero[07][07];
		diff_pixel[07][07][08] <= numero[07][08] > 7 ? numero[07][08] - 7 : 7 - numero[07][08];
		diff_pixel[07][07][09] <= numero[07][09] > 0 ? numero[07][09] - 0 : 0 - numero[07][09];
		diff_pixel[07][07][10] <= numero[07][10] > 0 ? numero[07][10] - 0 : 0 - numero[07][10];
		//diff_pixel[07][08][00] <= numero[08][00] > 11 ? numero[08][00] - 11 : 11 - numero[08][00];
		//diff_pixel[07][08][01] <= numero[08][01] > 12 ? numero[08][01] - 12 : 12 - numero[08][01];
		//diff_pixel[07][08][02] <= numero[08][02] > 45 ? numero[08][02] - 45 : 45 - numero[08][02];
		//diff_pixel[07][08][03] <= numero[08][03] > 99 ? numero[08][03] - 99 : 99 - numero[08][03];
		//diff_pixel[07][08][04] <= numero[08][04] > 130 ? numero[08][04] - 130 : 130 - numero[08][04];
		//diff_pixel[07][08][05] <= numero[08][05] > 128 ? numero[08][05] - 128 : 128 - numero[08][05];
		//diff_pixel[07][08][06] <= numero[08][06] > 94 ? numero[08][06] - 94 : 94 - numero[08][06];
		//diff_pixel[07][08][07] <= numero[08][07] > 43 ? numero[08][07] - 43 : 43 - numero[08][07];
		//diff_pixel[07][08][08] <= numero[08][08] > 8 ? numero[08][08] - 8 : 8 - numero[08][08];
		//diff_pixel[07][08][09] <= numero[08][09] > 0 ? numero[08][09] - 0 : 0 - numero[08][09];
		//diff_pixel[07][08][10] <= numero[08][10] > 0 ? numero[08][10] - 0 : 0 - numero[08][10];
		//diff_pixel[07][09][00] <= numero[09][00] > 0 ? numero[09][00] - 0 : 0 - numero[09][00];
		//diff_pixel[07][09][01] <= numero[09][01] > 14 ? numero[09][01] - 14 : 14 - numero[09][01];
		//diff_pixel[07][09][02] <= numero[09][02] > 49 ? numero[09][02] - 49 : 49 - numero[09][02];
		//diff_pixel[07][09][03] <= numero[09][03] > 101 ? numero[09][03] - 101 : 101 - numero[09][03];
		//diff_pixel[07][09][04] <= numero[09][04] > 130 ? numero[09][04] - 130 : 130 - numero[09][04];
		//diff_pixel[07][09][05] <= numero[09][05] > 128 ? numero[09][05] - 128 : 128 - numero[09][05];
		//diff_pixel[07][09][06] <= numero[09][06] > 92 ? numero[09][06] - 92 : 92 - numero[09][06];
		//diff_pixel[07][09][07] <= numero[09][07] > 40 ? numero[09][07] - 40 : 40 - numero[09][07];
		//diff_pixel[07][09][08] <= numero[09][08] > 7 ? numero[09][08] - 7 : 7 - numero[09][08];
		//diff_pixel[07][09][09] <= numero[09][09] > 0 ? numero[09][09] - 0 : 0 - numero[09][09];
		//diff_pixel[07][09][10] <= numero[09][10] > 0 ? numero[09][10] - 0 : 0 - numero[09][10];
		//diff_pixel[07][10][00] <= numero[10][00] > 0 ? numero[10][00] - 0 : 0 - numero[10][00];
		//diff_pixel[07][10][01] <= numero[10][01] > 2 ? numero[10][01] - 2 : 2 - numero[10][01];
		//diff_pixel[07][10][02] <= numero[10][02] > 28 ? numero[10][02] - 28 : 28 - numero[10][02];
		//diff_pixel[07][10][03] <= numero[10][03] > 63 ? numero[10][03] - 63 : 63 - numero[10][03];
		//diff_pixel[07][10][04] <= numero[10][04] > 85 ? numero[10][04] - 85 : 85 - numero[10][04];
		//diff_pixel[07][10][05] <= numero[10][05] > 85 ? numero[10][05] - 85 : 85 - numero[10][05];
		//diff_pixel[07][10][06] <= numero[10][06] > 60 ? numero[10][06] - 60 : 60 - numero[10][06];
		//diff_pixel[07][10][07] <= numero[10][07] > 24 ? numero[10][07] - 24 : 24 - numero[10][07];
		//diff_pixel[07][10][08] <= numero[10][08] > 2 ? numero[10][08] - 2 : 2 - numero[10][08];
		//diff_pixel[07][10][09] <= numero[10][09] > 0 ? numero[10][09] - 0 : 0 - numero[10][09];
//		
		//diff_pixel[08][00][00] <= numero[00][00] > 46 ? numero[00][00] - 46 : 46 - numero[00][00];
		//diff_pixel[08][00][01] <= numero[00][01] > 62 ? numero[00][01] - 62 : 62 - numero[00][01];
		//diff_pixel[08][00][02] <= numero[00][02] > 82 ? numero[00][02] - 82 : 82 - numero[00][02];
		//diff_pixel[08][00][03] <= numero[00][03] > 104 ? numero[00][03] - 104 : 104 - numero[00][03];
		//diff_pixel[08][00][04] <= numero[00][04] > 104 ? numero[00][04] - 104 : 104 - numero[00][04];
		//diff_pixel[08][00][05] <= numero[00][05] > 101 ? numero[00][05] - 101 : 101 - numero[00][05];
		//diff_pixel[08][00][06] <= numero[00][06] > 81 ? numero[00][06] - 81 : 81 - numero[00][06];
		//diff_pixel[08][00][07] <= numero[00][07] > 59 ? numero[00][07] - 59 : 59 - numero[00][07];
		//diff_pixel[08][00][08] <= numero[00][08] > 26 ? numero[00][08] - 26 : 26 - numero[00][08];
		//diff_pixel[08][00][09] <= numero[00][09] > 4 ? numero[00][09] - 4 : 4 - numero[00][09];
		//diff_pixel[08][00][10] <= numero[00][10] > 0 ? numero[00][10] - 0 : 0 - numero[00][10];
		//diff_pixel[08][01][00] <= numero[01][00] > 73 ? numero[01][00] - 73 : 73 - numero[01][00];
		//diff_pixel[08][01][01] <= numero[01][01] > 94 ? numero[01][01] - 94 : 94 - numero[01][01];
		//diff_pixel[08][01][02] <= numero[01][02] > 126 ? numero[01][02] - 126 : 126 - numero[01][02];
		//diff_pixel[08][01][03] <= numero[01][03] > 145 ? numero[01][03] - 145 : 145 - numero[01][03];
		//diff_pixel[08][01][04] <= numero[01][04] > 144 ? numero[01][04] - 144 : 144 - numero[01][04];
		//diff_pixel[08][01][05] <= numero[01][05] > 134 ? numero[01][05] - 134 : 134 - numero[01][05];
		//diff_pixel[08][01][06] <= numero[01][06] > 114 ? numero[01][06] - 114 : 114 - numero[01][06];
		//diff_pixel[08][01][07] <= numero[01][07] > 93 ? numero[01][07] - 93 : 93 - numero[01][07];
		//diff_pixel[08][01][08] <= numero[01][08] > 60 ? numero[01][08] - 60 : 60 - numero[01][08];
		//diff_pixel[08][01][09] <= numero[01][09] > 27 ? numero[01][09] - 27 : 27 - numero[01][09];
		//diff_pixel[08][01][10] <= numero[01][10] > 3 ? numero[01][10] - 3 : 3 - numero[01][10];
		diff_pixel[08][02][00] <= numero[02][00] > 117 ? numero[02][00] - 117 : 117 - numero[02][00];
		diff_pixel[08][02][01] <= numero[02][01] > 121 ? numero[02][01] - 121 : 121 - numero[02][01];
		diff_pixel[08][02][02] <= numero[02][02] > 114 ? numero[02][02] - 114 : 114 - numero[02][02];
		diff_pixel[08][02][03] <= numero[02][03] > 80 ? numero[02][03] - 80 : 80 - numero[02][03];
		diff_pixel[08][02][04] <= numero[02][04] > 36 ? numero[02][04] - 36 : 36 - numero[02][04];
		diff_pixel[08][02][05] <= numero[02][05] > 15 ? numero[02][05] - 15 : 15 - numero[02][05];
		diff_pixel[08][02][06] <= numero[02][06] > 27 ? numero[02][06] - 27 : 27 - numero[02][06];
		diff_pixel[08][02][07] <= numero[02][07] > 47 ? numero[02][07] - 47 : 47 - numero[02][07];
		diff_pixel[08][02][08] <= numero[02][08] > 70 ? numero[02][08] - 70 : 70 - numero[02][08];
		diff_pixel[08][02][09] <= numero[02][09] > 62 ? numero[02][09] - 62 : 62 - numero[02][09];
		diff_pixel[08][02][10] <= numero[02][10] > 36 ? numero[02][10] - 36 : 36 - numero[02][10];
		diff_pixel[08][03][00] <= numero[03][00] > 117 ? numero[03][00] - 117 : 117 - numero[03][00];
		diff_pixel[08][03][01] <= numero[03][01] > 149 ? numero[03][01] - 149 : 149 - numero[03][01];
		diff_pixel[08][03][02] <= numero[03][02] > 150 ? numero[03][02] - 150 : 150 - numero[03][02];
		diff_pixel[08][03][03] <= numero[03][03] > 124 ? numero[03][03] - 124 : 124 - numero[03][03];
		diff_pixel[08][03][04] <= numero[03][04] > 73 ? numero[03][04] - 73 : 73 - numero[03][04];
		diff_pixel[08][03][05] <= numero[03][05] > 35 ? numero[03][05] - 35 : 35 - numero[03][05];
		diff_pixel[08][03][06] <= numero[03][06] > 32 ? numero[03][06] - 32 : 32 - numero[03][06];
		diff_pixel[08][03][07] <= numero[03][07] > 43 ? numero[03][07] - 43 : 43 - numero[03][07];
		diff_pixel[08][03][08] <= numero[03][08] > 63 ? numero[03][08] - 63 : 63 - numero[03][08];
		diff_pixel[08][03][09] <= numero[03][09] > 59 ? numero[03][09] - 59 : 59 - numero[03][09];
		diff_pixel[08][03][10] <= numero[03][10] > 41 ? numero[03][10] - 41 : 41 - numero[03][10];
		diff_pixel[08][04][00] <= numero[04][00] > 77 ? numero[04][00] - 77 : 77 - numero[04][00];
		diff_pixel[08][04][01] <= numero[04][01] > 124 ? numero[04][01] - 124 : 124 - numero[04][01];
		diff_pixel[08][04][02] <= numero[04][02] > 151 ? numero[04][02] - 151 : 151 - numero[04][02];
		diff_pixel[08][04][03] <= numero[04][03] > 149 ? numero[04][03] - 149 : 149 - numero[04][03];
		diff_pixel[08][04][04] <= numero[04][04] > 125 ? numero[04][04] - 125 : 125 - numero[04][04];
		diff_pixel[08][04][05] <= numero[04][05] > 92 ? numero[04][05] - 92 : 92 - numero[04][05];
		diff_pixel[08][04][06] <= numero[04][06] > 77 ? numero[04][06] - 77 : 77 - numero[04][06];
		diff_pixel[08][04][07] <= numero[04][07] > 69 ? numero[04][07] - 69 : 69 - numero[04][07];
		diff_pixel[08][04][08] <= numero[04][08] > 70 ? numero[04][08] - 70 : 70 - numero[04][08];
		diff_pixel[08][04][09] <= numero[04][09] > 55 ? numero[04][09] - 55 : 55 - numero[04][09];
		diff_pixel[08][04][10] <= numero[04][10] > 41 ? numero[04][10] - 41 : 41 - numero[04][10];
		diff_pixel[08][05][00] <= numero[05][00] > 38 ? numero[05][00] - 38 : 38 - numero[05][00];
		diff_pixel[08][05][01] <= numero[05][01] > 82 ? numero[05][01] - 82 : 82 - numero[05][01];
		diff_pixel[08][05][02] <= numero[05][02] > 131 ? numero[05][02] - 131 : 131 - numero[05][02];
		diff_pixel[08][05][03] <= numero[05][03] > 162 ? numero[05][03] - 162 : 162 - numero[05][03];
		diff_pixel[08][05][04] <= numero[05][04] > 175 ? numero[05][04] - 175 : 175 - numero[05][04];
		diff_pixel[08][05][05] <= numero[05][05] > 170 ? numero[05][05] - 170 : 170 - numero[05][05];
		diff_pixel[08][05][06] <= numero[05][06] > 139 ? numero[05][06] - 139 : 139 - numero[05][06];
		diff_pixel[08][05][07] <= numero[05][07] > 105 ? numero[05][07] - 105 : 105 - numero[05][07];
		diff_pixel[08][05][08] <= numero[05][08] > 56 ? numero[05][08] - 56 : 56 - numero[05][08];
		diff_pixel[08][05][09] <= numero[05][09] > 15 ? numero[05][09] - 15 : 15 - numero[05][09];
		diff_pixel[08][05][10] <= numero[05][10] > 7 ? numero[05][10] - 7 : 7 - numero[05][10];
		diff_pixel[08][06][00] <= numero[06][00] > 51 ? numero[06][00] - 51 : 51 - numero[06][00];
		diff_pixel[08][06][01] <= numero[06][01] > 65 ? numero[06][01] - 65 : 65 - numero[06][01];
		diff_pixel[08][06][02] <= numero[06][02] > 73 ? numero[06][02] - 73 : 73 - numero[06][02];
		diff_pixel[08][06][03] <= numero[06][03] > 85 ? numero[06][03] - 85 : 85 - numero[06][03];
		diff_pixel[08][06][04] <= numero[06][04] > 105 ? numero[06][04] - 105 : 105 - numero[06][04];
		diff_pixel[08][06][05] <= numero[06][05] > 134 ? numero[06][05] - 134 : 134 - numero[06][05];
		diff_pixel[08][06][06] <= numero[06][06] > 154 ? numero[06][06] - 154 : 154 - numero[06][06];
		diff_pixel[08][06][07] <= numero[06][07] > 153 ? numero[06][07] - 153 : 153 - numero[06][07];
		diff_pixel[08][06][08] <= numero[06][08] > 138 ? numero[06][08] - 138 : 138 - numero[06][08];
		diff_pixel[08][06][09] <= numero[06][09] > 104 ? numero[06][09] - 104 : 104 - numero[06][09];
		diff_pixel[08][06][10] <= numero[06][10] > 85 ? numero[06][10] - 85 : 85 - numero[06][10];
		diff_pixel[08][07][00] <= numero[07][00] > 69 ? numero[07][00] - 69 : 69 - numero[07][00];
		diff_pixel[08][07][01] <= numero[07][01] > 64 ? numero[07][01] - 64 : 64 - numero[07][01];
		diff_pixel[08][07][02] <= numero[07][02] > 40 ? numero[07][02] - 40 : 40 - numero[07][02];
		diff_pixel[08][07][03] <= numero[07][03] > 32 ? numero[07][03] - 32 : 32 - numero[07][03];
		diff_pixel[08][07][04] <= numero[07][04] > 33 ? numero[07][04] - 33 : 33 - numero[07][04];
		diff_pixel[08][07][05] <= numero[07][05] > 68 ? numero[07][05] - 68 : 68 - numero[07][05];
		diff_pixel[08][07][06] <= numero[07][06] > 110 ? numero[07][06] - 110 : 110 - numero[07][06];
		diff_pixel[08][07][07] <= numero[07][07] > 138 ? numero[07][07] - 138 : 138 - numero[07][07];
		diff_pixel[08][07][08] <= numero[07][08] > 155 ? numero[07][08] - 155 : 155 - numero[07][08];
		diff_pixel[08][07][09] <= numero[07][09] > 141 ? numero[07][09] - 141 : 141 - numero[07][09];
		diff_pixel[08][07][10] <= numero[07][10] > 123 ? numero[07][10] - 123 : 123 - numero[07][10];
		//diff_pixel[08][08][00] <= numero[08][00] > 71 ? numero[08][00] - 71 : 71 - numero[08][00];
		//diff_pixel[08][08][01] <= numero[08][01] > 67 ? numero[08][01] - 67 : 67 - numero[08][01];
		//diff_pixel[08][08][02] <= numero[08][02] > 40 ? numero[08][02] - 40 : 40 - numero[08][02];
		//diff_pixel[08][08][03] <= numero[08][03] > 13 ? numero[08][03] - 13 : 13 - numero[08][03];
		//diff_pixel[08][08][04] <= numero[08][04] > 0 ? numero[08][04] - 0 : 0 - numero[08][04];
		//diff_pixel[08][08][05] <= numero[08][05] > 0 ? numero[08][05] - 0 : 0 - numero[08][05];
		//diff_pixel[08][08][06] <= numero[08][06] > 23 ? numero[08][06] - 23 : 23 - numero[08][06];
		//diff_pixel[08][08][07] <= numero[08][07] > 62 ? numero[08][07] - 62 : 62 - numero[08][07];
		//diff_pixel[08][08][08] <= numero[08][08] > 109 ? numero[08][08] - 109 : 109 - numero[08][08];
		//diff_pixel[08][08][09] <= numero[08][09] > 125 ? numero[08][09] - 125 : 125 - numero[08][09];
		//diff_pixel[08][08][10] <= numero[08][10] > 113 ? numero[08][10] - 113 : 113 - numero[08][10];
		//diff_pixel[08][09][00] <= numero[09][00] > 41 ? numero[09][00] - 41 : 41 - numero[09][00];
		//diff_pixel[08][09][01] <= numero[09][01] > 70 ? numero[09][01] - 70 : 70 - numero[09][01];
		//diff_pixel[08][09][02] <= numero[09][02] > 94 ? numero[09][02] - 94 : 94 - numero[09][02];
		//diff_pixel[08][09][03] <= numero[09][03] > 110 ? numero[09][03] - 110 : 110 - numero[09][03];
		//diff_pixel[08][09][04] <= numero[09][04] > 110 ? numero[09][04] - 110 : 110 - numero[09][04];
		//diff_pixel[08][09][05] <= numero[09][05] > 113 ? numero[09][05] - 113 : 113 - numero[09][05];
		//diff_pixel[08][09][06] <= numero[09][06] > 125 ? numero[09][06] - 125 : 125 - numero[09][06];
		//diff_pixel[08][09][07] <= numero[09][07] > 127 ? numero[09][07] - 127 : 127 - numero[09][07];
		//diff_pixel[08][09][08] <= numero[09][08] > 127 ? numero[09][08] - 127 : 127 - numero[09][08];
		//diff_pixel[08][09][09] <= numero[09][09] > 102 ? numero[09][09] - 102 : 102 - numero[09][09];
		//diff_pixel[08][09][10] <= numero[09][10] > 66 ? numero[09][10] - 66 : 66 - numero[09][10];
		//diff_pixel[08][10][00] <= numero[10][00] > 21 ? numero[10][00] - 21 : 21 - numero[10][00];
		//diff_pixel[08][10][01] <= numero[10][01] > 52 ? numero[10][01] - 52 : 52 - numero[10][01];
		//diff_pixel[08][10][02] <= numero[10][02] > 92 ? numero[10][02] - 92 : 92 - numero[10][02];
		//diff_pixel[08][10][03] <= numero[10][03] > 116 ? numero[10][03] - 116 : 116 - numero[10][03];
		//diff_pixel[08][10][04] <= numero[10][04] > 133 ? numero[10][04] - 133 : 133 - numero[10][04];
		//diff_pixel[08][10][05] <= numero[10][05] > 135 ? numero[10][05] - 135 : 135 - numero[10][05];
		//diff_pixel[08][10][06] <= numero[10][06] > 128 ? numero[10][06] - 128 : 128 - numero[10][06];
		//diff_pixel[08][10][07] <= numero[10][07] > 117 ? numero[10][07] - 117 : 117 - numero[10][07];
		//diff_pixel[08][10][08] <= numero[10][08] > 95 ? numero[10][08] - 95 : 95 - numero[10][08];
		//diff_pixel[08][10][09] <= numero[10][09] > 65 ? numero[10][09] - 65 : 65 - numero[10][09];
		//diff_pixel[08][10][10] <= numero[10][10] > 26 ? numero[10][10] - 26 : 26 - numero[10][10];
		
		//diff_pixel[09][00][00] <= numero[00][00] > 14 ? numero[00][00] - 14 : 14 - numero[00][00];
		//diff_pixel[09][00][01] <= numero[00][01] > 40 ? numero[00][01] - 40 : 40 - numero[00][01];
		//diff_pixel[09][00][02] <= numero[00][02] > 71 ? numero[00][02] - 71 : 71 - numero[00][02];
		//diff_pixel[09][00][03] <= numero[00][03] > 91 ? numero[00][03] - 91 : 91 - numero[00][03];
		//diff_pixel[09][00][04] <= numero[00][04] > 101 ? numero[00][04] - 101 : 101 - numero[00][04];
		//diff_pixel[09][00][05] <= numero[00][05] > 104 ? numero[00][05] - 104 : 104 - numero[00][05];
		//diff_pixel[09][00][06] <= numero[00][06] > 99 ? numero[00][06] - 99 : 99 - numero[00][06];
		//diff_pixel[09][00][07] <= numero[00][07] > 91 ? numero[00][07] - 91 : 91 - numero[00][07];
		//diff_pixel[09][00][08] <= numero[00][08] > 76 ? numero[00][08] - 76 : 76 - numero[00][08];
		//diff_pixel[09][00][09] <= numero[00][09] > 51 ? numero[00][09] - 51 : 51 - numero[00][09];
		//diff_pixel[09][00][10] <= numero[00][10] > 23 ? numero[00][10] - 23 : 23 - numero[00][10];
		//diff_pixel[09][01][00] <= numero[01][00] > 56 ? numero[01][00] - 56 : 56 - numero[01][00];
		//diff_pixel[09][01][01] <= numero[01][01] > 95 ? numero[01][01] - 95 : 95 - numero[01][01];
		//diff_pixel[09][01][02] <= numero[01][02] > 132 ? numero[01][02] - 132 : 132 - numero[01][02];
		//diff_pixel[09][01][03] <= numero[01][03] > 148 ? numero[01][03] - 148 : 148 - numero[01][03];
		//diff_pixel[09][01][04] <= numero[01][04] > 148 ? numero[01][04] - 148 : 148 - numero[01][04];
		//diff_pixel[09][01][05] <= numero[01][05] > 143 ? numero[01][05] - 143 : 143 - numero[01][05];
		//diff_pixel[09][01][06] <= numero[01][06] > 145 ? numero[01][06] - 145 : 145 - numero[01][06];
		//diff_pixel[09][01][07] <= numero[01][07] > 142 ? numero[01][07] - 142 : 142 - numero[01][07];
		//diff_pixel[09][01][08] <= numero[01][08] > 133 ? numero[01][08] - 133 : 133 - numero[01][08];
		//diff_pixel[09][01][09] <= numero[01][09] > 104 ? numero[01][09] - 104 : 104 - numero[01][09];
		//diff_pixel[09][01][10] <= numero[01][10] > 61 ? numero[01][10] - 61 : 61 - numero[01][10];
		diff_pixel[09][02][00] <= numero[02][00] > 97 ? numero[02][00] - 97 : 97 - numero[02][00];
		diff_pixel[09][02][01] <= numero[02][01] > 124 ? numero[02][01] - 124 : 124 - numero[02][01];
		diff_pixel[09][02][02] <= numero[02][02] > 123 ? numero[02][02] - 123 : 123 - numero[02][02];
		diff_pixel[09][02][03] <= numero[02][03] > 86 ? numero[02][03] - 86 : 86 - numero[02][03];
		diff_pixel[09][02][04] <= numero[02][04] > 44 ? numero[02][04] - 44 : 44 - numero[02][04];
		diff_pixel[09][02][05] <= numero[02][05] > 24 ? numero[02][05] - 24 : 24 - numero[02][05];
		diff_pixel[09][02][06] <= numero[02][06] > 33 ? numero[02][06] - 33 : 33 - numero[02][06];
		diff_pixel[09][02][07] <= numero[02][07] > 69 ? numero[02][07] - 69 : 69 - numero[02][07];
		diff_pixel[09][02][08] <= numero[02][08] > 112 ? numero[02][08] - 112 : 112 - numero[02][08];
		diff_pixel[09][02][09] <= numero[02][09] > 125 ? numero[02][09] - 125 : 125 - numero[02][09];
		diff_pixel[09][02][10] <= numero[02][10] > 107 ? numero[02][10] - 107 : 107 - numero[02][10];
		diff_pixel[09][03][00] <= numero[03][00] > 119 ? numero[03][00] - 119 : 119 - numero[03][00];
		diff_pixel[09][03][01] <= numero[03][01] > 130 ? numero[03][01] - 130 : 130 - numero[03][01];
		diff_pixel[09][03][02] <= numero[03][02] > 123 ? numero[03][02] - 123 : 123 - numero[03][02];
		diff_pixel[09][03][03] <= numero[03][03] > 83 ? numero[03][03] - 83 : 83 - numero[03][03];
		diff_pixel[09][03][04] <= numero[03][04] > 36 ? numero[03][04] - 36 : 36 - numero[03][04];
		diff_pixel[09][03][05] <= numero[03][05] > 12 ? numero[03][05] - 12 : 12 - numero[03][05];
		diff_pixel[09][03][06] <= numero[03][06] > 25 ? numero[03][06] - 25 : 25 - numero[03][06];
		diff_pixel[09][03][07] <= numero[03][07] > 65 ? numero[03][07] - 65 : 65 - numero[03][07];
		diff_pixel[09][03][08] <= numero[03][08] > 112 ? numero[03][08] - 112 : 112 - numero[03][08];
		diff_pixel[09][03][09] <= numero[03][09] > 129 ? numero[03][09] - 129 : 129 - numero[03][09];
		diff_pixel[09][03][10] <= numero[03][10] > 122 ? numero[03][10] - 122 : 122 - numero[03][10];
		diff_pixel[09][04][00] <= numero[04][00] > 92 ? numero[04][00] - 92 : 92 - numero[04][00];
		diff_pixel[09][04][01] <= numero[04][01] > 103 ? numero[04][01] - 103 : 103 - numero[04][01];
		diff_pixel[09][04][02] <= numero[04][02] > 116 ? numero[04][02] - 116 : 116 - numero[04][02];
		diff_pixel[09][04][03] <= numero[04][03] > 103 ? numero[04][03] - 103 : 103 - numero[04][03];
		diff_pixel[09][04][04] <= numero[04][04] > 77 ? numero[04][04] - 77 : 77 - numero[04][04];
		diff_pixel[09][04][05] <= numero[04][05] > 62 ? numero[04][05] - 62 : 62 - numero[04][05];
		diff_pixel[09][04][06] <= numero[04][06] > 68 ? numero[04][06] - 68 : 68 - numero[04][06];
		diff_pixel[09][04][07] <= numero[04][07] > 95 ? numero[04][07] - 95 : 95 - numero[04][07];
		diff_pixel[09][04][08] <= numero[04][08] > 126 ? numero[04][08] - 126 : 126 - numero[04][08];
		diff_pixel[09][04][09] <= numero[04][09] > 130 ? numero[04][09] - 130 : 130 - numero[04][09];
		diff_pixel[09][04][10] <= numero[04][10] > 121 ? numero[04][10] - 121 : 121 - numero[04][10];
		diff_pixel[09][05][00] <= numero[05][00] > 51 ? numero[05][00] - 51 : 51 - numero[05][00];
		diff_pixel[09][05][01] <= numero[05][01] > 76 ? numero[05][01] - 76 : 76 - numero[05][01];
		diff_pixel[09][05][02] <= numero[05][02] > 125 ? numero[05][02] - 125 : 125 - numero[05][02];
		diff_pixel[09][05][03] <= numero[05][03] > 159 ? numero[05][03] - 159 : 159 - numero[05][03];
		diff_pixel[09][05][04] <= numero[05][04] > 175 ? numero[05][04] - 175 : 175 - numero[05][04];
		diff_pixel[09][05][05] <= numero[05][05] > 175 ? numero[05][05] - 175 : 175 - numero[05][05];
		diff_pixel[09][05][06] <= numero[05][06] > 170 ? numero[05][06] - 170 : 170 - numero[05][06];
		diff_pixel[09][05][07] <= numero[05][07] > 174 ? numero[05][07] - 174 : 174 - numero[05][07];
		diff_pixel[09][05][08] <= numero[05][08] > 172 ? numero[05][08] - 172 : 172 - numero[05][08];
		diff_pixel[09][05][09] <= numero[05][09] > 151 ? numero[05][09] - 151 : 151 - numero[05][09];
		diff_pixel[09][05][10] <= numero[05][10] > 128 ? numero[05][10] - 128 : 128 - numero[05][10];
		diff_pixel[09][06][00] <= numero[06][00] > 19 ? numero[06][00] - 19 : 19 - numero[06][00];
		diff_pixel[09][06][01] <= numero[06][01] > 19 ? numero[06][01] - 19 : 19 - numero[06][01];
		diff_pixel[09][06][02] <= numero[06][02] > 39 ? numero[06][02] - 39 : 39 - numero[06][02];
		diff_pixel[09][06][03] <= numero[06][03] > 56 ? numero[06][03] - 56 : 56 - numero[06][03];
		diff_pixel[09][06][04] <= numero[06][04] > 63 ? numero[06][04] - 63 : 63 - numero[06][04];
		diff_pixel[09][06][05] <= numero[06][05] > 66 ? numero[06][05] - 66 : 66 - numero[06][05];
		diff_pixel[09][06][06] <= numero[06][06] > 81 ? numero[06][06] - 81 : 81 - numero[06][06];
		diff_pixel[09][06][07] <= numero[06][07] > 104 ? numero[06][07] - 104 : 104 - numero[06][07];
		diff_pixel[09][06][08] <= numero[06][08] > 133 ? numero[06][08] - 133 : 133 - numero[06][08];
		diff_pixel[09][06][09] <= numero[06][09] > 135 ? numero[06][09] - 135 : 135 - numero[06][09];
		diff_pixel[09][06][10] <= numero[06][10] > 126 ? numero[06][10] - 126 : 126 - numero[06][10];
		diff_pixel[09][07][00] <= numero[07][00] > 0 ? numero[07][00] - 0 : 0 - numero[07][00];
		diff_pixel[09][07][01] <= numero[07][01] > 0 ? numero[07][01] - 0 : 0 - numero[07][01];
		diff_pixel[09][07][02] <= numero[07][02] > 0 ? numero[07][02] - 0 : 0 - numero[07][02];
		diff_pixel[09][07][03] <= numero[07][03] > 0 ? numero[07][03] - 0 : 0 - numero[07][03];
		diff_pixel[09][07][04] <= numero[07][04] > 0 ? numero[07][04] - 0 : 0 - numero[07][04];
		diff_pixel[09][07][05] <= numero[07][05] > 10 ? numero[07][05] - 10 : 10 - numero[07][05];
		diff_pixel[09][07][06] <= numero[07][06] > 41 ? numero[07][06] - 41 : 41 - numero[07][06];
		diff_pixel[09][07][07] <= numero[07][07] > 79 ? numero[07][07] - 79 : 79 - numero[07][07];
		diff_pixel[09][07][08] <= numero[07][08] > 114 ? numero[07][08] - 114 : 114 - numero[07][08];
		diff_pixel[09][07][09] <= numero[07][09] > 116 ? numero[07][09] - 116 : 116 - numero[07][09];
		diff_pixel[09][07][10] <= numero[07][10] > 100 ? numero[07][10] - 100 : 100 - numero[07][10];
		//diff_pixel[09][08][00] <= numero[08][00] > 0 ? numero[08][00] - 0 : 0 - numero[08][00];
		//diff_pixel[09][08][01] <= numero[08][01] > 0 ? numero[08][01] - 0 : 0 - numero[08][01];
		//diff_pixel[09][08][02] <= numero[08][02] > 0 ? numero[08][02] - 0 : 0 - numero[08][02];
		//diff_pixel[09][08][03] <= numero[08][03] > 0 ? numero[08][03] - 0 : 0 - numero[08][03];
		//diff_pixel[09][08][04] <= numero[08][04] > 13 ? numero[08][04] - 13 : 13 - numero[08][04];
		//diff_pixel[09][08][05] <= numero[08][05] > 42 ? numero[08][05] - 42 : 42 - numero[08][05];
		//diff_pixel[09][08][06] <= numero[08][06] > 93 ? numero[08][06] - 93 : 93 - numero[08][06];
		//diff_pixel[09][08][07] <= numero[08][07] > 129 ? numero[08][07] - 129 : 129 - numero[08][07];
		//diff_pixel[09][08][08] <= numero[08][08] > 136 ? numero[08][08] - 136 : 136 - numero[08][08];
		//diff_pixel[09][08][09] <= numero[08][09] > 107 ? numero[08][09] - 107 : 107 - numero[08][09];
		//diff_pixel[09][08][10] <= numero[08][10] > 51 ? numero[08][10] - 51 : 51 - numero[08][10];
		//diff_pixel[09][09][00] <= numero[09][00] > 16 ? numero[09][00] - 16 : 16 - numero[09][00];
		//diff_pixel[09][09][01] <= numero[09][01] > 49 ? numero[09][01] - 49 : 49 - numero[09][01];
		//diff_pixel[09][09][02] <= numero[09][02] > 87 ? numero[09][02] - 87 : 87 - numero[09][02];
		//diff_pixel[09][09][03] <= numero[09][03] > 111 ? numero[09][03] - 111 : 111 - numero[09][03];
		//diff_pixel[09][09][04] <= numero[09][04] > 131 ? numero[09][04] - 131 : 131 - numero[09][04];
		//diff_pixel[09][09][05] <= numero[09][05] > 138 ? numero[09][05] - 138 : 138 - numero[09][05];
		//diff_pixel[09][09][06] <= numero[09][06] > 134 ? numero[09][06] - 134 : 134 - numero[09][06];
		//diff_pixel[09][09][07] <= numero[09][07] > 119 ? numero[09][07] - 119 : 119 - numero[09][07];
		//diff_pixel[09][09][08] <= numero[09][08] > 87 ? numero[09][08] - 87 : 87 - numero[09][08];
		//diff_pixel[09][09][09] <= numero[09][09] > 50 ? numero[09][09] - 50 : 50 - numero[09][09];
		//diff_pixel[09][09][10] <= numero[09][10] > 15 ? numero[09][10] - 15 : 15 - numero[09][10];
		//diff_pixel[09][10][00] <= numero[10][00] > 20 ? numero[10][00] - 20 : 20 - numero[10][00];
		//diff_pixel[09][10][01] <= numero[10][01] > 51 ? numero[10][01] - 51 : 51 - numero[10][01];
		//diff_pixel[09][10][02] <= numero[10][02] > 85 ? numero[10][02] - 85 : 85 - numero[10][02];
		//diff_pixel[09][10][03] <= numero[10][03] > 110 ? numero[10][03] - 110 : 110 - numero[10][03];
		//diff_pixel[09][10][04] <= numero[10][04] > 122 ? numero[10][04] - 122 : 122 - numero[10][04];
		//diff_pixel[09][10][05] <= numero[10][05] > 121 ? numero[10][05] - 121 : 121 - numero[10][05];
		//diff_pixel[09][10][06] <= numero[10][06] > 101 ? numero[10][06] - 101 : 101 - numero[10][06];
		//diff_pixel[09][10][07] <= numero[10][07] > 75 ? numero[10][07] - 75 : 75 - numero[10][07];
		//diff_pixel[09][10][08] <= numero[10][08] > 39 ? numero[10][08] - 39 : 39 - numero[10][08];
		//diff_pixel[09][10][09] <= numero[10][09] > 11 ? numero[10][09] - 11 : 11 - numero[10][09];
		//diff_pixel[09][10][10] <= numero[10][10] > 0 ? numero[10][10] - 0 : 0 - numero[10][10];
		
	end
	
endmodule
