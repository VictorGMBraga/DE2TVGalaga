module Diferenca6(
	input  [7:0] numero[3:1][10:0][10:0],
	output [15:0] diff_pixel[3:1][10:0][10:0]
	);
	
	DiferencaEuclidiana diferencaEuclidiana_1_0_0(numero[1][0][0],19,diff_pixel[1][0][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_1(numero[1][0][1],30,diff_pixel[1][0][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_2(numero[1][0][2],41,diff_pixel[1][0][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_3(numero[1][0][3],69,diff_pixel[1][0][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_4(numero[1][0][4],84,diff_pixel[1][0][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_5(numero[1][0][5],100,diff_pixel[1][0][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_6(numero[1][0][6],104,diff_pixel[1][0][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_7(numero[1][0][7],96,diff_pixel[1][0][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_8(numero[1][0][8],73,diff_pixel[1][0][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_9(numero[1][0][9],48,diff_pixel[1][0][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_10(numero[1][0][10],21,diff_pixel[1][0][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_0(numero[1][1][0],9,diff_pixel[1][1][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_1(numero[1][1][1],35,diff_pixel[1][1][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_2(numero[1][1][2],70,diff_pixel[1][1][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_3(numero[1][1][3],111,diff_pixel[1][1][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_4(numero[1][1][4],136,diff_pixel[1][1][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_5(numero[1][1][5],143,diff_pixel[1][1][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_6(numero[1][1][6],142,diff_pixel[1][1][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_7(numero[1][1][7],125,diff_pixel[1][1][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_8(numero[1][1][8],102,diff_pixel[1][1][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_9(numero[1][1][9],70,diff_pixel[1][1][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_10(numero[1][1][10],32,diff_pixel[1][1][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_0(numero[1][2][0],44,diff_pixel[1][2][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_1(numero[1][2][1],72,diff_pixel[1][2][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_2(numero[1][2][2],111,diff_pixel[1][2][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_3(numero[1][2][3],126,diff_pixel[1][2][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_4(numero[1][2][4],106,diff_pixel[1][2][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_5(numero[1][2][5],59,diff_pixel[1][2][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_6(numero[1][2][6],23,diff_pixel[1][2][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_7(numero[1][2][7],2,diff_pixel[1][2][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_8(numero[1][2][8],0,diff_pixel[1][2][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_9(numero[1][2][9],0,diff_pixel[1][2][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_10(numero[1][2][10],0,diff_pixel[1][2][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_0(numero[1][3][0],100,diff_pixel[1][3][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_1(numero[1][3][1],111,diff_pixel[1][3][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_2(numero[1][3][2],120,diff_pixel[1][3][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_3(numero[1][3][3],100,diff_pixel[1][3][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_4(numero[1][3][4],59,diff_pixel[1][3][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_5(numero[1][3][5],21,diff_pixel[1][3][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_6(numero[1][3][6],0,diff_pixel[1][3][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_7(numero[1][3][7],0,diff_pixel[1][3][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_8(numero[1][3][8],0,diff_pixel[1][3][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_9(numero[1][3][9],0,diff_pixel[1][3][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_10(numero[1][3][10],0,diff_pixel[1][3][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_0(numero[1][4][0],119,diff_pixel[1][4][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_1(numero[1][4][1],129,diff_pixel[1][4][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_2(numero[1][4][2],129,diff_pixel[1][4][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_3(numero[1][4][3],107,diff_pixel[1][4][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_4(numero[1][4][4],73,diff_pixel[1][4][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_5(numero[1][4][5],53,diff_pixel[1][4][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_6(numero[1][4][6],45,diff_pixel[1][4][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_7(numero[1][4][7],43,diff_pixel[1][4][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_8(numero[1][4][8],36,diff_pixel[1][4][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_9(numero[1][4][9],21,diff_pixel[1][4][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_10(numero[1][4][10],15,diff_pixel[1][4][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_0(numero[1][5][0],126,diff_pixel[1][5][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_1(numero[1][5][1],148,diff_pixel[1][5][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_2(numero[1][5][2],170,diff_pixel[1][5][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_3(numero[1][5][3],179,diff_pixel[1][5][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_4(numero[1][5][4],174,diff_pixel[1][5][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_5(numero[1][5][5],168,diff_pixel[1][5][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_6(numero[1][5][6],168,diff_pixel[1][5][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_7(numero[1][5][7],157,diff_pixel[1][5][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_8(numero[1][5][8],129,diff_pixel[1][5][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_9(numero[1][5][9],86,diff_pixel[1][5][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_10(numero[1][5][10],48,diff_pixel[1][5][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_0(numero[1][6][0],122,diff_pixel[1][6][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_1(numero[1][6][1],134,diff_pixel[1][6][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_2(numero[1][6][2],136,diff_pixel[1][6][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_3(numero[1][6][3],117,diff_pixel[1][6][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_4(numero[1][6][4],86,diff_pixel[1][6][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_5(numero[1][6][5],71,diff_pixel[1][6][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_6(numero[1][6][6],81,diff_pixel[1][6][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_7(numero[1][6][7],101,diff_pixel[1][6][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_8(numero[1][6][8],124,diff_pixel[1][6][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_9(numero[1][6][9],117,diff_pixel[1][6][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_10(numero[1][6][10],99,diff_pixel[1][6][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_0(numero[1][7][0],115,diff_pixel[1][7][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_1(numero[1][7][1],126,diff_pixel[1][7][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_2(numero[1][7][2],118,diff_pixel[1][7][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_3(numero[1][7][3],80,diff_pixel[1][7][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_4(numero[1][7][4],33,diff_pixel[1][7][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_5(numero[1][7][5],9,diff_pixel[1][7][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_6(numero[1][7][6],20,diff_pixel[1][7][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_7(numero[1][7][7],60,diff_pixel[1][7][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_8(numero[1][7][8],108,diff_pixel[1][7][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_9(numero[1][7][9],125,diff_pixel[1][7][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_10(numero[1][7][10],119,diff_pixel[1][7][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_0(numero[1][8][0],105,diff_pixel[1][8][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_1(numero[1][8][1],131,diff_pixel[1][8][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_2(numero[1][8][2],120,diff_pixel[1][8][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_3(numero[1][8][3],78,diff_pixel[1][8][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_4(numero[1][8][4],28,diff_pixel[1][8][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_5(numero[1][8][5],4,diff_pixel[1][8][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_6(numero[1][8][6],22,diff_pixel[1][8][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_7(numero[1][8][7],62,diff_pixel[1][8][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_8(numero[1][8][8],115,diff_pixel[1][8][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_9(numero[1][8][9],134,diff_pixel[1][8][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_10(numero[1][8][10],118,diff_pixel[1][8][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_0(numero[1][9][0],58,diff_pixel[1][9][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_1(numero[1][9][1],95,diff_pixel[1][9][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_2(numero[1][9][2],131,diff_pixel[1][9][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_3(numero[1][9][3],142,diff_pixel[1][9][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_4(numero[1][9][4],138,diff_pixel[1][9][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_5(numero[1][9][5],134,diff_pixel[1][9][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_6(numero[1][9][6],134,diff_pixel[1][9][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_7(numero[1][9][7],136,diff_pixel[1][9][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_8(numero[1][9][8],134,diff_pixel[1][9][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_9(numero[1][9][9],110,diff_pixel[1][9][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_10(numero[1][9][10],66,diff_pixel[1][9][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_0(numero[1][10][0],16,diff_pixel[1][10][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_1(numero[1][10][1],47,diff_pixel[1][10][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_2(numero[1][10][2],80,diff_pixel[1][10][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_3(numero[1][10][3],103,diff_pixel[1][10][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_4(numero[1][10][4],113,diff_pixel[1][10][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_5(numero[1][10][5],115,diff_pixel[1][10][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_6(numero[1][10][6],119,diff_pixel[1][10][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_7(numero[1][10][7],108,diff_pixel[1][10][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_8(numero[1][10][8],95,diff_pixel[1][10][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_9(numero[1][10][9],64,diff_pixel[1][10][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_10(numero[1][10][10],30,diff_pixel[1][10][10]);

	DiferencaEuclidiana diferencaEuclidiana_2_0_0(numero[2][0][0],0,diff_pixel[2][0][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_1(numero[2][0][1],0,diff_pixel[2][0][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_2(numero[2][0][2],16,diff_pixel[2][0][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_3(numero[2][0][3],44,diff_pixel[2][0][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_4(numero[2][0][4],73,diff_pixel[2][0][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_5(numero[2][0][5],89,diff_pixel[2][0][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_6(numero[2][0][6],100,diff_pixel[2][0][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_7(numero[2][0][7],92,diff_pixel[2][0][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_8(numero[2][0][8],77,diff_pixel[2][0][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_9(numero[2][0][9],52,diff_pixel[2][0][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_10(numero[2][0][10],22,diff_pixel[2][0][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_0(numero[2][1][0],3,diff_pixel[2][1][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_1(numero[2][1][1],29,diff_pixel[2][1][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_2(numero[2][1][2],66,diff_pixel[2][1][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_3(numero[2][1][3],107,diff_pixel[2][1][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_4(numero[2][1][4],135,diff_pixel[2][1][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_5(numero[2][1][5],142,diff_pixel[2][1][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_6(numero[2][1][6],142,diff_pixel[2][1][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_7(numero[2][1][7],125,diff_pixel[2][1][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_8(numero[2][1][8],103,diff_pixel[2][1][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_9(numero[2][1][9],71,diff_pixel[2][1][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_10(numero[2][1][10],32,diff_pixel[2][1][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_0(numero[2][2][0],39,diff_pixel[2][2][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_1(numero[2][2][1],67,diff_pixel[2][2][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_2(numero[2][2][2],110,diff_pixel[2][2][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_3(numero[2][2][3],125,diff_pixel[2][2][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_4(numero[2][2][4],109,diff_pixel[2][2][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_5(numero[2][2][5],62,diff_pixel[2][2][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_6(numero[2][2][6],23,diff_pixel[2][2][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_7(numero[2][2][7],2,diff_pixel[2][2][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_8(numero[2][2][8],0,diff_pixel[2][2][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_9(numero[2][2][9],0,diff_pixel[2][2][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_10(numero[2][2][10],0,diff_pixel[2][2][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_0(numero[2][3][0],91,diff_pixel[2][3][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_1(numero[2][3][1],102,diff_pixel[2][3][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_2(numero[2][3][2],113,diff_pixel[2][3][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_3(numero[2][3][3],93,diff_pixel[2][3][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_4(numero[2][3][4],57,diff_pixel[2][3][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_5(numero[2][3][5],19,diff_pixel[2][3][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_6(numero[2][3][6],0,diff_pixel[2][3][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_7(numero[2][3][7],0,diff_pixel[2][3][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_8(numero[2][3][8],0,diff_pixel[2][3][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_9(numero[2][3][9],0,diff_pixel[2][3][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_10(numero[2][3][10],0,diff_pixel[2][3][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_0(numero[2][4][0],124,diff_pixel[2][4][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_1(numero[2][4][1],134,diff_pixel[2][4][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_2(numero[2][4][2],135,diff_pixel[2][4][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_3(numero[2][4][3],113,diff_pixel[2][4][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_4(numero[2][4][4],79,diff_pixel[2][4][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_5(numero[2][4][5],59,diff_pixel[2][4][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_6(numero[2][4][6],49,diff_pixel[2][4][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_7(numero[2][4][7],47,diff_pixel[2][4][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_8(numero[2][4][8],40,diff_pixel[2][4][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_9(numero[2][4][9],25,diff_pixel[2][4][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_10(numero[2][4][10],21,diff_pixel[2][4][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_0(numero[2][5][0],125,diff_pixel[2][5][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_1(numero[2][5][1],147,diff_pixel[2][5][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_2(numero[2][5][2],169,diff_pixel[2][5][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_3(numero[2][5][3],178,diff_pixel[2][5][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_4(numero[2][5][4],174,diff_pixel[2][5][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_5(numero[2][5][5],168,diff_pixel[2][5][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_6(numero[2][5][6],169,diff_pixel[2][5][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_7(numero[2][5][7],158,diff_pixel[2][5][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_8(numero[2][5][8],133,diff_pixel[2][5][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_9(numero[2][5][9],90,diff_pixel[2][5][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_10(numero[2][5][10],52,diff_pixel[2][5][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_0(numero[2][6][0],123,diff_pixel[2][6][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_1(numero[2][6][1],135,diff_pixel[2][6][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_2(numero[2][6][2],136,diff_pixel[2][6][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_3(numero[2][6][3],117,diff_pixel[2][6][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_4(numero[2][6][4],86,diff_pixel[2][6][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_5(numero[2][6][5],71,diff_pixel[2][6][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_6(numero[2][6][6],80,diff_pixel[2][6][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_7(numero[2][6][7],100,diff_pixel[2][6][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_8(numero[2][6][8],120,diff_pixel[2][6][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_9(numero[2][6][9],113,diff_pixel[2][6][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_10(numero[2][6][10],98,diff_pixel[2][6][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_0(numero[2][7][0],116,diff_pixel[2][7][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_1(numero[2][7][1],127,diff_pixel[2][7][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_2(numero[2][7][2],117,diff_pixel[2][7][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_3(numero[2][7][3],79,diff_pixel[2][7][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_4(numero[2][7][4],29,diff_pixel[2][7][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_5(numero[2][7][5],5,diff_pixel[2][7][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_6(numero[2][7][6],19,diff_pixel[2][7][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_7(numero[2][7][7],59,diff_pixel[2][7][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_8(numero[2][7][8],108,diff_pixel[2][7][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_9(numero[2][7][9],125,diff_pixel[2][7][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_10(numero[2][7][10],123,diff_pixel[2][7][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_0(numero[2][8][0],100,diff_pixel[2][8][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_1(numero[2][8][1],126,diff_pixel[2][8][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_2(numero[2][8][2],119,diff_pixel[2][8][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_3(numero[2][8][3],77,diff_pixel[2][8][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_4(numero[2][8][4],29,diff_pixel[2][8][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_5(numero[2][8][5],5,diff_pixel[2][8][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_6(numero[2][8][6],18,diff_pixel[2][8][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_7(numero[2][8][7],58,diff_pixel[2][8][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_8(numero[2][8][8],107,diff_pixel[2][8][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_9(numero[2][8][9],126,diff_pixel[2][8][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_10(numero[2][8][10],112,diff_pixel[2][8][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_0(numero[2][9][0],53,diff_pixel[2][9][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_1(numero[2][9][1],90,diff_pixel[2][9][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_2(numero[2][9][2],122,diff_pixel[2][9][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_3(numero[2][9][3],133,diff_pixel[2][9][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_4(numero[2][9][4],129,diff_pixel[2][9][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_5(numero[2][9][5],125,diff_pixel[2][9][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_6(numero[2][9][6],128,diff_pixel[2][9][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_7(numero[2][9][7],130,diff_pixel[2][9][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_8(numero[2][9][8],129,diff_pixel[2][9][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_9(numero[2][9][9],105,diff_pixel[2][9][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_10(numero[2][9][10],65,diff_pixel[2][9][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_0(numero[2][10][0],18,diff_pixel[2][10][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_1(numero[2][10][1],49,diff_pixel[2][10][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_2(numero[2][10][2],88,diff_pixel[2][10][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_3(numero[2][10][3],111,diff_pixel[2][10][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_4(numero[2][10][4],126,diff_pixel[2][10][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_5(numero[2][10][5],128,diff_pixel[2][10][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_6(numero[2][10][6],126,diff_pixel[2][10][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_7(numero[2][10][7],115,diff_pixel[2][10][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_8(numero[2][10][8],97,diff_pixel[2][10][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_9(numero[2][10][9],66,diff_pixel[2][10][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_10(numero[2][10][10],26,diff_pixel[2][10][10]);

	DiferencaEuclidiana diferencaEuclidiana_3_0_0(numero[3][0][0],0,diff_pixel[3][0][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_1(numero[3][0][1],0,diff_pixel[3][0][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_2(numero[3][0][2],22,diff_pixel[3][0][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_3(numero[3][0][3],50,diff_pixel[3][0][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_4(numero[3][0][4],81,diff_pixel[3][0][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_5(numero[3][0][5],97,diff_pixel[3][0][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_6(numero[3][0][6],105,diff_pixel[3][0][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_7(numero[3][0][7],97,diff_pixel[3][0][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_8(numero[3][0][8],78,diff_pixel[3][0][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_9(numero[3][0][9],53,diff_pixel[3][0][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_10(numero[3][0][10],22,diff_pixel[3][0][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_0(numero[3][1][0],5,diff_pixel[3][1][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_1(numero[3][1][1],31,diff_pixel[3][1][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_2(numero[3][1][2],69,diff_pixel[3][1][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_3(numero[3][1][3],110,diff_pixel[3][1][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_4(numero[3][1][4],139,diff_pixel[3][1][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_5(numero[3][1][5],146,diff_pixel[3][1][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_6(numero[3][1][6],146,diff_pixel[3][1][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_7(numero[3][1][7],129,diff_pixel[3][1][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_8(numero[3][1][8],105,diff_pixel[3][1][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_9(numero[3][1][9],73,diff_pixel[3][1][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_10(numero[3][1][10],34,diff_pixel[3][1][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_0(numero[3][2][0],51,diff_pixel[3][2][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_1(numero[3][2][1],79,diff_pixel[3][2][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_2(numero[3][2][2],119,diff_pixel[3][2][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_3(numero[3][2][3],134,diff_pixel[3][2][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_4(numero[3][2][4],115,diff_pixel[3][2][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_5(numero[3][2][5],68,diff_pixel[3][2][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_6(numero[3][2][6],30,diff_pixel[3][2][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_7(numero[3][2][7],9,diff_pixel[3][2][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_8(numero[3][2][8],2,diff_pixel[3][2][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_9(numero[3][2][9],3,diff_pixel[3][2][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_10(numero[3][2][10],0,diff_pixel[3][2][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_0(numero[3][3][0],98,diff_pixel[3][3][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_1(numero[3][3][1],109,diff_pixel[3][3][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_2(numero[3][3][2],124,diff_pixel[3][3][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_3(numero[3][3][3],104,diff_pixel[3][3][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_4(numero[3][3][4],68,diff_pixel[3][3][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_5(numero[3][3][5],30,diff_pixel[3][3][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_6(numero[3][3][6],7,diff_pixel[3][3][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_7(numero[3][3][7],0,diff_pixel[3][3][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_8(numero[3][3][8],0,diff_pixel[3][3][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_9(numero[3][3][9],0,diff_pixel[3][3][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_10(numero[3][3][10],4,diff_pixel[3][3][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_0(numero[3][4][0],131,diff_pixel[3][4][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_1(numero[3][4][1],141,diff_pixel[3][4][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_2(numero[3][4][2],137,diff_pixel[3][4][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_3(numero[3][4][3],115,diff_pixel[3][4][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_4(numero[3][4][4],75,diff_pixel[3][4][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_5(numero[3][4][5],55,diff_pixel[3][4][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_6(numero[3][4][6],48,diff_pixel[3][4][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_7(numero[3][4][7],46,diff_pixel[3][4][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_8(numero[3][4][8],41,diff_pixel[3][4][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_9(numero[3][4][9],26,diff_pixel[3][4][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_10(numero[3][4][10],17,diff_pixel[3][4][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_0(numero[3][5][0],125,diff_pixel[3][5][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_1(numero[3][5][1],147,diff_pixel[3][5][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_2(numero[3][5][2],171,diff_pixel[3][5][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_3(numero[3][5][3],180,diff_pixel[3][5][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_4(numero[3][5][4],178,diff_pixel[3][5][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_5(numero[3][5][5],172,diff_pixel[3][5][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_6(numero[3][5][6],173,diff_pixel[3][5][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_7(numero[3][5][7],162,diff_pixel[3][5][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_8(numero[3][5][8],136,diff_pixel[3][5][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_9(numero[3][5][9],93,diff_pixel[3][5][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_10(numero[3][5][10],51,diff_pixel[3][5][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_0(numero[3][6][0],123,diff_pixel[3][6][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_1(numero[3][6][1],135,diff_pixel[3][6][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_2(numero[3][6][2],134,diff_pixel[3][6][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_3(numero[3][6][3],115,diff_pixel[3][6][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_4(numero[3][6][4],82,diff_pixel[3][6][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_5(numero[3][6][5],67,diff_pixel[3][6][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_6(numero[3][6][6],80,diff_pixel[3][6][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_7(numero[3][6][7],100,diff_pixel[3][6][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_8(numero[3][6][8],123,diff_pixel[3][6][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_9(numero[3][6][9],116,diff_pixel[3][6][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_10(numero[3][6][10],102,diff_pixel[3][6][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_0(numero[3][7][0],107,diff_pixel[3][7][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_1(numero[3][7][1],118,diff_pixel[3][7][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_2(numero[3][7][2],113,diff_pixel[3][7][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_3(numero[3][7][3],75,diff_pixel[3][7][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_4(numero[3][7][4],30,diff_pixel[3][7][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_5(numero[3][7][5],6,diff_pixel[3][7][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_6(numero[3][7][6],23,diff_pixel[3][7][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_7(numero[3][7][7],63,diff_pixel[3][7][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_8(numero[3][7][8],117,diff_pixel[3][7][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_9(numero[3][7][9],134,diff_pixel[3][7][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_10(numero[3][7][10],126,diff_pixel[3][7][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_0(numero[3][8][0],110,diff_pixel[3][8][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_1(numero[3][8][1],136,diff_pixel[3][8][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_2(numero[3][8][2],123,diff_pixel[3][8][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_3(numero[3][8][3],81,diff_pixel[3][8][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_4(numero[3][8][4],27,diff_pixel[3][8][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_5(numero[3][8][5],3,diff_pixel[3][8][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_6(numero[3][8][6],15,diff_pixel[3][8][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_7(numero[3][8][7],55,diff_pixel[3][8][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_8(numero[3][8][8],103,diff_pixel[3][8][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_9(numero[3][8][9],122,diff_pixel[3][8][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_10(numero[3][8][10],118,diff_pixel[3][8][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_0(numero[3][9][0],48,diff_pixel[3][9][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_1(numero[3][9][1],85,diff_pixel[3][9][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_2(numero[3][9][2],123,diff_pixel[3][9][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_3(numero[3][9][3],134,diff_pixel[3][9][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_4(numero[3][9][4],132,diff_pixel[3][9][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_5(numero[3][9][5],128,diff_pixel[3][9][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_6(numero[3][9][6],134,diff_pixel[3][9][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_7(numero[3][9][7],136,diff_pixel[3][9][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_8(numero[3][9][8],139,diff_pixel[3][9][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_9(numero[3][9][9],115,diff_pixel[3][9][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_10(numero[3][9][10],74,diff_pixel[3][9][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_0(numero[3][10][0],33,diff_pixel[3][10][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_1(numero[3][10][1],64,diff_pixel[3][10][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_2(numero[3][10][2],92,diff_pixel[3][10][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_3(numero[3][10][3],115,diff_pixel[3][10][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_4(numero[3][10][4],120,diff_pixel[3][10][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_5(numero[3][10][5],122,diff_pixel[3][10][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_6(numero[3][10][6],115,diff_pixel[3][10][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_7(numero[3][10][7],104,diff_pixel[3][10][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_8(numero[3][10][8],81,diff_pixel[3][10][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_9(numero[3][10][9],50,diff_pixel[3][10][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_10(numero[3][10][10],23,diff_pixel[3][10][10]);
	

endmodule

