module Diferenca4(
	input  [7:0] numero[3:1][10:0][10:0],
	output [15:0] diff_pixel[3:1][10:0][10:0]
	);
	
	DiferencaEuclidiana diferencaEuclidiana_1_0_0(numero[1][0][0],14,diff_pixel[1][0][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_1(numero[1][0][1],14,diff_pixel[1][0][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_2(numero[1][0][2],10,diff_pixel[1][0][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_3(numero[1][0][3],24,diff_pixel[1][0][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_4(numero[1][0][4],40,diff_pixel[1][0][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_5(numero[1][0][5],70,diff_pixel[1][0][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_6(numero[1][0][6],89,diff_pixel[1][0][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_7(numero[1][0][7],91,diff_pixel[1][0][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_8(numero[1][0][8],78,diff_pixel[1][0][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_9(numero[1][0][9],50,diff_pixel[1][0][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_0_10(numero[1][0][10],19,diff_pixel[1][0][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_0(numero[1][1][0],0,diff_pixel[1][1][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_1(numero[1][1][1],0,diff_pixel[1][1][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_2(numero[1][1][2],12,diff_pixel[1][1][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_3(numero[1][1][3],46,diff_pixel[1][1][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_4(numero[1][1][4],86,diff_pixel[1][1][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_5(numero[1][1][5],134,diff_pixel[1][1][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_6(numero[1][1][6],166,diff_pixel[1][1][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_7(numero[1][1][7],167,diff_pixel[1][1][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_8(numero[1][1][8],143,diff_pixel[1][1][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_9(numero[1][1][9],95,diff_pixel[1][1][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_1_10(numero[1][1][10],44,diff_pixel[1][1][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_0(numero[1][2][0],0,diff_pixel[1][2][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_1(numero[1][2][1],20,diff_pixel[1][2][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_2(numero[1][2][2],49,diff_pixel[1][2][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_3(numero[1][2][3],98,diff_pixel[1][2][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_4(numero[1][2][4],139,diff_pixel[1][2][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_5(numero[1][2][5],168,diff_pixel[1][2][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_6(numero[1][2][6],182,diff_pixel[1][2][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_7(numero[1][2][7],168,diff_pixel[1][2][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_8(numero[1][2][8],136,diff_pixel[1][2][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_9(numero[1][2][9],91,diff_pixel[1][2][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_2_10(numero[1][2][10],44,diff_pixel[1][2][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_0(numero[1][3][0],24,diff_pixel[1][3][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_1(numero[1][3][1],51,diff_pixel[1][3][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_2(numero[1][3][2],91,diff_pixel[1][3][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_3(numero[1][3][3],117,diff_pixel[1][3][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_4(numero[1][3][4],132,diff_pixel[1][3][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_5(numero[1][3][5],127,diff_pixel[1][3][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_6(numero[1][3][6],136,diff_pixel[1][3][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_7(numero[1][3][7],139,diff_pixel[1][3][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_8(numero[1][3][8],126,diff_pixel[1][3][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_9(numero[1][3][9],93,diff_pixel[1][3][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_3_10(numero[1][3][10],51,diff_pixel[1][3][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_0(numero[1][4][0],78,diff_pixel[1][4][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_1(numero[1][4][1],98,diff_pixel[1][4][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_2(numero[1][4][2],116,diff_pixel[1][4][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_3(numero[1][4][3],112,diff_pixel[1][4][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_4(numero[1][4][4],92,diff_pixel[1][4][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_5(numero[1][4][5],77,diff_pixel[1][4][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_6(numero[1][4][6],99,diff_pixel[1][4][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_7(numero[1][4][7],120,diff_pixel[1][4][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_8(numero[1][4][8],126,diff_pixel[1][4][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_9(numero[1][4][9],97,diff_pixel[1][4][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_4_10(numero[1][4][10],63,diff_pixel[1][4][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_0(numero[1][5][0],123,diff_pixel[1][5][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_1(numero[1][5][1],128,diff_pixel[1][5][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_2(numero[1][5][2],119,diff_pixel[1][5][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_3(numero[1][5][3],84,diff_pixel[1][5][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_4(numero[1][5][4],52,diff_pixel[1][5][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_5(numero[1][5][5],51,diff_pixel[1][5][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_6(numero[1][5][6],86,diff_pixel[1][5][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_7(numero[1][5][7],123,diff_pixel[1][5][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_8(numero[1][5][8],128,diff_pixel[1][5][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_9(numero[1][5][9],97,diff_pixel[1][5][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_5_10(numero[1][5][10],59,diff_pixel[1][5][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_0(numero[1][6][0],121,diff_pixel[1][6][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_1(numero[1][6][1],137,diff_pixel[1][6][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_2(numero[1][6][2],147,diff_pixel[1][6][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_3(numero[1][6][3],140,diff_pixel[1][6][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_4(numero[1][6][4],124,diff_pixel[1][6][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_5(numero[1][6][5],122,diff_pixel[1][6][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_6(numero[1][6][6],140,diff_pixel[1][6][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_7(numero[1][6][7],155,diff_pixel[1][6][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_8(numero[1][6][8],157,diff_pixel[1][6][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_9(numero[1][6][9],130,diff_pixel[1][6][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_6_10(numero[1][6][10],103,diff_pixel[1][6][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_0(numero[1][7][0],84,diff_pixel[1][7][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_1(numero[1][7][1],103,diff_pixel[1][7][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_2(numero[1][7][2],116,diff_pixel[1][7][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_3(numero[1][7][3],124,diff_pixel[1][7][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_4(numero[1][7][4],124,diff_pixel[1][7][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_5(numero[1][7][5],131,diff_pixel[1][7][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_6(numero[1][7][6],150,diff_pixel[1][7][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_7(numero[1][7][7],161,diff_pixel[1][7][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_8(numero[1][7][8],161,diff_pixel[1][7][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_9(numero[1][7][9],135,diff_pixel[1][7][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_7_10(numero[1][7][10],106,diff_pixel[1][7][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_0(numero[1][8][0],0,diff_pixel[1][8][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_1(numero[1][8][1],0,diff_pixel[1][8][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_2(numero[1][8][2],0,diff_pixel[1][8][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_3(numero[1][8][3],0,diff_pixel[1][8][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_4(numero[1][8][4],4,diff_pixel[1][8][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_5(numero[1][8][5],33,diff_pixel[1][8][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_6(numero[1][8][6],83,diff_pixel[1][8][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_7(numero[1][8][7],118,diff_pixel[1][8][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_8(numero[1][8][8],122,diff_pixel[1][8][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_9(numero[1][8][9],91,diff_pixel[1][8][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_8_10(numero[1][8][10],43,diff_pixel[1][8][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_0(numero[1][9][0],0,diff_pixel[1][9][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_1(numero[1][9][1],0,diff_pixel[1][9][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_2(numero[1][9][2],0,diff_pixel[1][9][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_3(numero[1][9][3],0,diff_pixel[1][9][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_4(numero[1][9][4],3,diff_pixel[1][9][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_5(numero[1][9][5],31,diff_pixel[1][9][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_6(numero[1][9][6],83,diff_pixel[1][9][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_7(numero[1][9][7],119,diff_pixel[1][9][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_8(numero[1][9][8],126,diff_pixel[1][9][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_9(numero[1][9][9],97,diff_pixel[1][9][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_9_10(numero[1][9][10],48,diff_pixel[1][9][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_0(numero[1][10][0],0,diff_pixel[1][10][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_1(numero[1][10][1],0,diff_pixel[1][10][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_2(numero[1][10][2],0,diff_pixel[1][10][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_3(numero[1][10][3],0,diff_pixel[1][10][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_4(numero[1][10][4],4,diff_pixel[1][10][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_5(numero[1][10][5],24,diff_pixel[1][10][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_6(numero[1][10][6],58,diff_pixel[1][10][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_7(numero[1][10][7],82,diff_pixel[1][10][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_8(numero[1][10][8],83,diff_pixel[1][10][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_9(numero[1][10][9],62,diff_pixel[1][10][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_10_10(numero[1][10][10],29,diff_pixel[1][10][10]);

	DiferencaEuclidiana diferencaEuclidiana_2_0_0(numero[2][0][0],0,diff_pixel[2][0][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_1(numero[2][0][1],0,diff_pixel[2][0][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_2(numero[2][0][2],0,diff_pixel[2][0][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_3(numero[2][0][3],7,diff_pixel[2][0][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_4(numero[2][0][4],34,diff_pixel[2][0][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_5(numero[2][0][5],64,diff_pixel[2][0][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_6(numero[2][0][6],88,diff_pixel[2][0][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_7(numero[2][0][7],90,diff_pixel[2][0][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_8(numero[2][0][8],79,diff_pixel[2][0][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_9(numero[2][0][9],51,diff_pixel[2][0][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_0_10(numero[2][0][10],20,diff_pixel[2][0][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_0(numero[2][1][0],0,diff_pixel[2][1][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_1(numero[2][1][1],0,diff_pixel[2][1][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_2(numero[2][1][2],12,diff_pixel[2][1][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_3(numero[2][1][3],46,diff_pixel[2][1][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_4(numero[2][1][4],87,diff_pixel[2][1][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_5(numero[2][1][5],135,diff_pixel[2][1][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_6(numero[2][1][6],167,diff_pixel[2][1][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_7(numero[2][1][7],168,diff_pixel[2][1][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_8(numero[2][1][8],144,diff_pixel[2][1][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_9(numero[2][1][9],96,diff_pixel[2][1][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_1_10(numero[2][1][10],44,diff_pixel[2][1][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_0(numero[2][2][0],0,diff_pixel[2][2][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_1(numero[2][2][1],14,diff_pixel[2][2][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_2(numero[2][2][2],47,diff_pixel[2][2][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_3(numero[2][2][3],96,diff_pixel[2][2][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_4(numero[2][2][4],139,diff_pixel[2][2][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_5(numero[2][2][5],168,diff_pixel[2][2][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_6(numero[2][2][6],183,diff_pixel[2][2][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_7(numero[2][2][7],169,diff_pixel[2][2][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_8(numero[2][2][8],141,diff_pixel[2][2][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_9(numero[2][2][9],96,diff_pixel[2][2][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_2_10(numero[2][2][10],45,diff_pixel[2][2][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_0(numero[2][3][0],26,diff_pixel[2][3][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_1(numero[2][3][1],53,diff_pixel[2][3][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_2(numero[2][3][2],91,diff_pixel[2][3][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_3(numero[2][3][3],117,diff_pixel[2][3][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_4(numero[2][3][4],131,diff_pixel[2][3][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_5(numero[2][3][5],126,diff_pixel[2][3][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_6(numero[2][3][6],136,diff_pixel[2][3][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_7(numero[2][3][7],139,diff_pixel[2][3][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_8(numero[2][3][8],131,diff_pixel[2][3][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_9(numero[2][3][9],98,diff_pixel[2][3][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_3_10(numero[2][3][10],55,diff_pixel[2][3][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_0(numero[2][4][0],64,diff_pixel[2][4][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_1(numero[2][4][1],84,diff_pixel[2][4][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_2(numero[2][4][2],114,diff_pixel[2][4][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_3(numero[2][4][3],110,diff_pixel[2][4][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_4(numero[2][4][4],101,diff_pixel[2][4][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_5(numero[2][4][5],86,diff_pixel[2][4][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_6(numero[2][4][6],104,diff_pixel[2][4][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_7(numero[2][4][7],125,diff_pixel[2][4][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_8(numero[2][4][8],129,diff_pixel[2][4][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_9(numero[2][4][9],100,diff_pixel[2][4][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_4_10(numero[2][4][10],58,diff_pixel[2][4][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_0(numero[2][5][0],114,diff_pixel[2][5][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_1(numero[2][5][1],119,diff_pixel[2][5][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_2(numero[2][5][2],113,diff_pixel[2][5][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_3(numero[2][5][3],78,diff_pixel[2][5][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_4(numero[2][5][4],50,diff_pixel[2][5][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_5(numero[2][5][5],49,diff_pixel[2][5][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_6(numero[2][5][6],86,diff_pixel[2][5][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_7(numero[2][5][7],123,diff_pixel[2][5][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_8(numero[2][5][8],129,diff_pixel[2][5][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_9(numero[2][5][9],98,diff_pixel[2][5][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_5_10(numero[2][5][10],59,diff_pixel[2][5][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_0(numero[2][6][0],124,diff_pixel[2][6][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_1(numero[2][6][1],140,diff_pixel[2][6][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_2(numero[2][6][2],153,diff_pixel[2][6][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_3(numero[2][6][3],146,diff_pixel[2][6][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_4(numero[2][6][4],135,diff_pixel[2][6][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_5(numero[2][6][5],133,diff_pixel[2][6][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_6(numero[2][6][6],147,diff_pixel[2][6][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_7(numero[2][6][7],162,diff_pixel[2][6][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_8(numero[2][6][8],160,diff_pixel[2][6][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_9(numero[2][6][9],133,diff_pixel[2][6][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_6_10(numero[2][6][10],103,diff_pixel[2][6][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_0(numero[2][7][0],79,diff_pixel[2][7][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_1(numero[2][7][1],98,diff_pixel[2][7][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_2(numero[2][7][2],115,diff_pixel[2][7][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_3(numero[2][7][3],123,diff_pixel[2][7][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_4(numero[2][7][4],130,diff_pixel[2][7][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_5(numero[2][7][5],137,diff_pixel[2][7][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_6(numero[2][7][6],151,diff_pixel[2][7][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_7(numero[2][7][7],162,diff_pixel[2][7][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_8(numero[2][7][8],162,diff_pixel[2][7][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_9(numero[2][7][9],136,diff_pixel[2][7][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_7_10(numero[2][7][10],102,diff_pixel[2][7][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_0(numero[2][8][0],0,diff_pixel[2][8][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_1(numero[2][8][1],0,diff_pixel[2][8][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_2(numero[2][8][2],0,diff_pixel[2][8][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_3(numero[2][8][3],0,diff_pixel[2][8][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_4(numero[2][8][4],13,diff_pixel[2][8][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_5(numero[2][8][5],42,diff_pixel[2][8][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_6(numero[2][8][6],92,diff_pixel[2][8][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_7(numero[2][8][7],127,diff_pixel[2][8][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_8(numero[2][8][8],131,diff_pixel[2][8][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_9(numero[2][8][9],100,diff_pixel[2][8][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_8_10(numero[2][8][10],48,diff_pixel[2][8][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_0(numero[2][9][0],0,diff_pixel[2][9][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_1(numero[2][9][1],0,diff_pixel[2][9][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_2(numero[2][9][2],0,diff_pixel[2][9][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_3(numero[2][9][3],0,diff_pixel[2][9][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_4(numero[2][9][4],12,diff_pixel[2][9][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_5(numero[2][9][5],40,diff_pixel[2][9][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_6(numero[2][9][6],89,diff_pixel[2][9][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_7(numero[2][9][7],125,diff_pixel[2][9][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_8(numero[2][9][8],131,diff_pixel[2][9][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_9(numero[2][9][9],102,diff_pixel[2][9][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_9_10(numero[2][9][10],49,diff_pixel[2][9][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_0(numero[2][10][0],0,diff_pixel[2][10][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_1(numero[2][10][1],0,diff_pixel[2][10][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_2(numero[2][10][2],0,diff_pixel[2][10][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_3(numero[2][10][3],0,diff_pixel[2][10][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_4(numero[2][10][4],4,diff_pixel[2][10][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_5(numero[2][10][5],24,diff_pixel[2][10][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_6(numero[2][10][6],59,diff_pixel[2][10][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_7(numero[2][10][7],83,diff_pixel[2][10][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_8(numero[2][10][8],87,diff_pixel[2][10][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_9(numero[2][10][9],66,diff_pixel[2][10][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_10_10(numero[2][10][10],30,diff_pixel[2][10][10]);

	DiferencaEuclidiana diferencaEuclidiana_3_0_0(numero[3][0][0],0,diff_pixel[3][0][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_1(numero[3][0][1],0,diff_pixel[3][0][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_2(numero[3][0][2],0,diff_pixel[3][0][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_3(numero[3][0][3],6,diff_pixel[3][0][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_4(numero[3][0][4],32,diff_pixel[3][0][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_5(numero[3][0][5],62,diff_pixel[3][0][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_6(numero[3][0][6],86,diff_pixel[3][0][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_7(numero[3][0][7],88,diff_pixel[3][0][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_8(numero[3][0][8],79,diff_pixel[3][0][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_9(numero[3][0][9],51,diff_pixel[3][0][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_0_10(numero[3][0][10],20,diff_pixel[3][0][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_0(numero[3][1][0],0,diff_pixel[3][1][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_1(numero[3][1][1],0,diff_pixel[3][1][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_2(numero[3][1][2],10,diff_pixel[3][1][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_3(numero[3][1][3],44,diff_pixel[3][1][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_4(numero[3][1][4],85,diff_pixel[3][1][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_5(numero[3][1][5],133,diff_pixel[3][1][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_6(numero[3][1][6],167,diff_pixel[3][1][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_7(numero[3][1][7],168,diff_pixel[3][1][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_8(numero[3][1][8],144,diff_pixel[3][1][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_9(numero[3][1][9],96,diff_pixel[3][1][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_1_10(numero[3][1][10],44,diff_pixel[3][1][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_0(numero[3][2][0],0,diff_pixel[3][2][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_1(numero[3][2][1],20,diff_pixel[3][2][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_2(numero[3][2][2],54,diff_pixel[3][2][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_3(numero[3][2][3],103,diff_pixel[3][2][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_4(numero[3][2][4],146,diff_pixel[3][2][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_5(numero[3][2][5],175,diff_pixel[3][2][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_6(numero[3][2][6],183,diff_pixel[3][2][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_7(numero[3][2][7],169,diff_pixel[3][2][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_8(numero[3][2][8],131,diff_pixel[3][2][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_9(numero[3][2][9],86,diff_pixel[3][2][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_2_10(numero[3][2][10],38,diff_pixel[3][2][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_0(numero[3][3][0],15,diff_pixel[3][3][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_1(numero[3][3][1],42,diff_pixel[3][3][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_2(numero[3][3][2],87,diff_pixel[3][3][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_3(numero[3][3][3],113,diff_pixel[3][3][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_4(numero[3][3][4],133,diff_pixel[3][3][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_5(numero[3][3][5],128,diff_pixel[3][3][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_6(numero[3][3][6],143,diff_pixel[3][3][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_7(numero[3][3][7],146,diff_pixel[3][3][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_8(numero[3][3][8],138,diff_pixel[3][3][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_9(numero[3][3][9],105,diff_pixel[3][3][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_3_10(numero[3][3][10],56,diff_pixel[3][3][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_0(numero[3][4][0],87,diff_pixel[3][4][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_1(numero[3][4][1],107,diff_pixel[3][4][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_2(numero[3][4][2],125,diff_pixel[3][4][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_3(numero[3][4][3],121,diff_pixel[3][4][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_4(numero[3][4][4],102,diff_pixel[3][4][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_5(numero[3][4][5],87,diff_pixel[3][4][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_6(numero[3][4][6],94,diff_pixel[3][4][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_7(numero[3][4][7],115,diff_pixel[3][4][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_8(numero[3][4][8],106,diff_pixel[3][4][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_9(numero[3][4][9],77,diff_pixel[3][4][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_4_10(numero[3][4][10],49,diff_pixel[3][4][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_0(numero[3][5][0],115,diff_pixel[3][5][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_1(numero[3][5][1],120,diff_pixel[3][5][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_2(numero[3][5][2],119,diff_pixel[3][5][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_3(numero[3][5][3],84,diff_pixel[3][5][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_4(numero[3][5][4],59,diff_pixel[3][5][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_5(numero[3][5][5],58,diff_pixel[3][5][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_6(numero[3][5][6],90,diff_pixel[3][5][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_7(numero[3][5][7],127,diff_pixel[3][5][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_8(numero[3][5][8],129,diff_pixel[3][5][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_9(numero[3][5][9],98,diff_pixel[3][5][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_5_10(numero[3][5][10],59,diff_pixel[3][5][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_0(numero[3][6][0],134,diff_pixel[3][6][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_1(numero[3][6][1],150,diff_pixel[3][6][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_2(numero[3][6][2],155,diff_pixel[3][6][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_3(numero[3][6][3],148,diff_pixel[3][6][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_4(numero[3][6][4],127,diff_pixel[3][6][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_5(numero[3][6][5],125,diff_pixel[3][6][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_6(numero[3][6][6],136,diff_pixel[3][6][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_7(numero[3][6][7],151,diff_pixel[3][6][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_8(numero[3][6][8],146,diff_pixel[3][6][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_9(numero[3][6][9],119,diff_pixel[3][6][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_6_10(numero[3][6][10],96,diff_pixel[3][6][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_0(numero[3][7][0],89,diff_pixel[3][7][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_1(numero[3][7][1],108,diff_pixel[3][7][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_2(numero[3][7][2],122,diff_pixel[3][7][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_3(numero[3][7][3],130,diff_pixel[3][7][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_4(numero[3][7][4],132,diff_pixel[3][7][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_5(numero[3][7][5],139,diff_pixel[3][7][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_6(numero[3][7][6],149,diff_pixel[3][7][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_7(numero[3][7][7],160,diff_pixel[3][7][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_8(numero[3][7][8],153,diff_pixel[3][7][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_9(numero[3][7][9],127,diff_pixel[3][7][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_7_10(numero[3][7][10],101,diff_pixel[3][7][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_0(numero[3][8][0],0,diff_pixel[3][8][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_1(numero[3][8][1],0,diff_pixel[3][8][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_2(numero[3][8][2],0,diff_pixel[3][8][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_3(numero[3][8][3],0,diff_pixel[3][8][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_4(numero[3][8][4],10,diff_pixel[3][8][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_5(numero[3][8][5],39,diff_pixel[3][8][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_6(numero[3][8][6],89,diff_pixel[3][8][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_7(numero[3][8][7],124,diff_pixel[3][8][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_8(numero[3][8][8],126,diff_pixel[3][8][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_9(numero[3][8][9],95,diff_pixel[3][8][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_8_10(numero[3][8][10],38,diff_pixel[3][8][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_0(numero[3][9][0],0,diff_pixel[3][9][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_1(numero[3][9][1],0,diff_pixel[3][9][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_2(numero[3][9][2],0,diff_pixel[3][9][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_3(numero[3][9][3],0,diff_pixel[3][9][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_4(numero[3][9][4],9,diff_pixel[3][9][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_5(numero[3][9][5],37,diff_pixel[3][9][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_6(numero[3][9][6],83,diff_pixel[3][9][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_7(numero[3][9][7],119,diff_pixel[3][9][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_8(numero[3][9][8],119,diff_pixel[3][9][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_9(numero[3][9][9],90,diff_pixel[3][9][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_9_10(numero[3][9][10],40,diff_pixel[3][9][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_0(numero[3][10][0],0,diff_pixel[3][10][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_1(numero[3][10][1],0,diff_pixel[3][10][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_2(numero[3][10][2],0,diff_pixel[3][10][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_3(numero[3][10][3],0,diff_pixel[3][10][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_4(numero[3][10][4],6,diff_pixel[3][10][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_5(numero[3][10][5],26,diff_pixel[3][10][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_6(numero[3][10][6],63,diff_pixel[3][10][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_7(numero[3][10][7],87,diff_pixel[3][10][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_8(numero[3][10][8],90,diff_pixel[3][10][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_9(numero[3][10][9],69,diff_pixel[3][10][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_10_10(numero[3][10][10],28,diff_pixel[3][10][10]);
	

endmodule

