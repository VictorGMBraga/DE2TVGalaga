module checkNum(input [7:1]numero[7:1][3:1][10:0][10:0] );
endmodule