module Diferenca6(
	input  [7:0] numero[10:0][10:0],
	output [7:0] diff_pixel[10:0][10:0]
	);
	
	DiferencaEuclidiana diferencaEuclidiana_0_0(numero[0][0],19,diff_pixel[0][0]);
	DiferencaEuclidiana diferencaEuclidiana_0_1(numero[0][1],30,diff_pixel[0][1]);
	DiferencaEuclidiana diferencaEuclidiana_0_2(numero[0][2],41,diff_pixel[0][2]);
	DiferencaEuclidiana diferencaEuclidiana_0_3(numero[0][3],69,diff_pixel[0][3]);
	DiferencaEuclidiana diferencaEuclidiana_0_4(numero[0][4],84,diff_pixel[0][4]);
	DiferencaEuclidiana diferencaEuclidiana_0_5(numero[0][5],100,diff_pixel[0][5]);
	DiferencaEuclidiana diferencaEuclidiana_0_6(numero[0][6],104,diff_pixel[0][6]);
	DiferencaEuclidiana diferencaEuclidiana_0_7(numero[0][7],96,diff_pixel[0][7]);
	DiferencaEuclidiana diferencaEuclidiana_0_8(numero[0][8],73,diff_pixel[0][8]);
	DiferencaEuclidiana diferencaEuclidiana_0_9(numero[0][9],48,diff_pixel[0][9]);
	DiferencaEuclidiana diferencaEuclidiana_0_10(numero[0][10],21,diff_pixel[0][10]);
	DiferencaEuclidiana diferencaEuclidiana_1_0(numero[1][0],9,diff_pixel[1][0]);
	DiferencaEuclidiana diferencaEuclidiana_1_1(numero[1][1],35,diff_pixel[1][1]);
	DiferencaEuclidiana diferencaEuclidiana_1_2(numero[1][2],70,diff_pixel[1][2]);
	DiferencaEuclidiana diferencaEuclidiana_1_3(numero[1][3],111,diff_pixel[1][3]);
	DiferencaEuclidiana diferencaEuclidiana_1_4(numero[1][4],136,diff_pixel[1][4]);
	DiferencaEuclidiana diferencaEuclidiana_1_5(numero[1][5],143,diff_pixel[1][5]);
	DiferencaEuclidiana diferencaEuclidiana_1_6(numero[1][6],142,diff_pixel[1][6]);
	DiferencaEuclidiana diferencaEuclidiana_1_7(numero[1][7],125,diff_pixel[1][7]);
	DiferencaEuclidiana diferencaEuclidiana_1_8(numero[1][8],102,diff_pixel[1][8]);
	DiferencaEuclidiana diferencaEuclidiana_1_9(numero[1][9],70,diff_pixel[1][9]);
	DiferencaEuclidiana diferencaEuclidiana_1_10(numero[1][10],32,diff_pixel[1][10]);
	DiferencaEuclidiana diferencaEuclidiana_2_0(numero[2][0],44,diff_pixel[2][0]);
	DiferencaEuclidiana diferencaEuclidiana_2_1(numero[2][1],72,diff_pixel[2][1]);
	DiferencaEuclidiana diferencaEuclidiana_2_2(numero[2][2],111,diff_pixel[2][2]);
	DiferencaEuclidiana diferencaEuclidiana_2_3(numero[2][3],126,diff_pixel[2][3]);
	DiferencaEuclidiana diferencaEuclidiana_2_4(numero[2][4],106,diff_pixel[2][4]);
	DiferencaEuclidiana diferencaEuclidiana_2_5(numero[2][5],59,diff_pixel[2][5]);
	DiferencaEuclidiana diferencaEuclidiana_2_6(numero[2][6],23,diff_pixel[2][6]);
	DiferencaEuclidiana diferencaEuclidiana_2_7(numero[2][7],2,diff_pixel[2][7]);
	DiferencaEuclidiana diferencaEuclidiana_2_8(numero[2][8],0,diff_pixel[2][8]);
	DiferencaEuclidiana diferencaEuclidiana_2_9(numero[2][9],0,diff_pixel[2][9]);
	DiferencaEuclidiana diferencaEuclidiana_2_10(numero[2][10],0,diff_pixel[2][10]);
	DiferencaEuclidiana diferencaEuclidiana_3_0(numero[3][0],100,diff_pixel[3][0]);
	DiferencaEuclidiana diferencaEuclidiana_3_1(numero[3][1],111,diff_pixel[3][1]);
	DiferencaEuclidiana diferencaEuclidiana_3_2(numero[3][2],120,diff_pixel[3][2]);
	DiferencaEuclidiana diferencaEuclidiana_3_3(numero[3][3],100,diff_pixel[3][3]);
	DiferencaEuclidiana diferencaEuclidiana_3_4(numero[3][4],59,diff_pixel[3][4]);
	DiferencaEuclidiana diferencaEuclidiana_3_5(numero[3][5],21,diff_pixel[3][5]);
	DiferencaEuclidiana diferencaEuclidiana_3_6(numero[3][6],0,diff_pixel[3][6]);
	DiferencaEuclidiana diferencaEuclidiana_3_7(numero[3][7],0,diff_pixel[3][7]);
	DiferencaEuclidiana diferencaEuclidiana_3_8(numero[3][8],0,diff_pixel[3][8]);
	DiferencaEuclidiana diferencaEuclidiana_3_9(numero[3][9],0,diff_pixel[3][9]);
	DiferencaEuclidiana diferencaEuclidiana_3_10(numero[3][10],0,diff_pixel[3][10]);
	DiferencaEuclidiana diferencaEuclidiana_4_0(numero[4][0],119,diff_pixel[4][0]);
	DiferencaEuclidiana diferencaEuclidiana_4_1(numero[4][1],129,diff_pixel[4][1]);
	DiferencaEuclidiana diferencaEuclidiana_4_2(numero[4][2],129,diff_pixel[4][2]);
	DiferencaEuclidiana diferencaEuclidiana_4_3(numero[4][3],107,diff_pixel[4][3]);
	DiferencaEuclidiana diferencaEuclidiana_4_4(numero[4][4],73,diff_pixel[4][4]);
	DiferencaEuclidiana diferencaEuclidiana_4_5(numero[4][5],53,diff_pixel[4][5]);
	DiferencaEuclidiana diferencaEuclidiana_4_6(numero[4][6],45,diff_pixel[4][6]);
	DiferencaEuclidiana diferencaEuclidiana_4_7(numero[4][7],43,diff_pixel[4][7]);
	DiferencaEuclidiana diferencaEuclidiana_4_8(numero[4][8],36,diff_pixel[4][8]);
	DiferencaEuclidiana diferencaEuclidiana_4_9(numero[4][9],21,diff_pixel[4][9]);
	DiferencaEuclidiana diferencaEuclidiana_4_10(numero[4][10],15,diff_pixel[4][10]);
	DiferencaEuclidiana diferencaEuclidiana_5_0(numero[5][0],126,diff_pixel[5][0]);
	DiferencaEuclidiana diferencaEuclidiana_5_1(numero[5][1],148,diff_pixel[5][1]);
	DiferencaEuclidiana diferencaEuclidiana_5_2(numero[5][2],170,diff_pixel[5][2]);
	DiferencaEuclidiana diferencaEuclidiana_5_3(numero[5][3],179,diff_pixel[5][3]);
	DiferencaEuclidiana diferencaEuclidiana_5_4(numero[5][4],174,diff_pixel[5][4]);
	DiferencaEuclidiana diferencaEuclidiana_5_5(numero[5][5],168,diff_pixel[5][5]);
	DiferencaEuclidiana diferencaEuclidiana_5_6(numero[5][6],168,diff_pixel[5][6]);
	DiferencaEuclidiana diferencaEuclidiana_5_7(numero[5][7],157,diff_pixel[5][7]);
	DiferencaEuclidiana diferencaEuclidiana_5_8(numero[5][8],129,diff_pixel[5][8]);
	DiferencaEuclidiana diferencaEuclidiana_5_9(numero[5][9],86,diff_pixel[5][9]);
	DiferencaEuclidiana diferencaEuclidiana_5_10(numero[5][10],48,diff_pixel[5][10]);
	DiferencaEuclidiana diferencaEuclidiana_6_0(numero[6][0],122,diff_pixel[6][0]);
	DiferencaEuclidiana diferencaEuclidiana_6_1(numero[6][1],134,diff_pixel[6][1]);
	DiferencaEuclidiana diferencaEuclidiana_6_2(numero[6][2],136,diff_pixel[6][2]);
	DiferencaEuclidiana diferencaEuclidiana_6_3(numero[6][3],117,diff_pixel[6][3]);
	DiferencaEuclidiana diferencaEuclidiana_6_4(numero[6][4],86,diff_pixel[6][4]);
	DiferencaEuclidiana diferencaEuclidiana_6_5(numero[6][5],71,diff_pixel[6][5]);
	DiferencaEuclidiana diferencaEuclidiana_6_6(numero[6][6],81,diff_pixel[6][6]);
	DiferencaEuclidiana diferencaEuclidiana_6_7(numero[6][7],101,diff_pixel[6][7]);
	DiferencaEuclidiana diferencaEuclidiana_6_8(numero[6][8],124,diff_pixel[6][8]);
	DiferencaEuclidiana diferencaEuclidiana_6_9(numero[6][9],117,diff_pixel[6][9]);
	DiferencaEuclidiana diferencaEuclidiana_6_10(numero[6][10],99,diff_pixel[6][10]);
	DiferencaEuclidiana diferencaEuclidiana_7_0(numero[7][0],115,diff_pixel[7][0]);
	DiferencaEuclidiana diferencaEuclidiana_7_1(numero[7][1],126,diff_pixel[7][1]);
	DiferencaEuclidiana diferencaEuclidiana_7_2(numero[7][2],118,diff_pixel[7][2]);
	DiferencaEuclidiana diferencaEuclidiana_7_3(numero[7][3],80,diff_pixel[7][3]);
	DiferencaEuclidiana diferencaEuclidiana_7_4(numero[7][4],33,diff_pixel[7][4]);
	DiferencaEuclidiana diferencaEuclidiana_7_5(numero[7][5],9,diff_pixel[7][5]);
	DiferencaEuclidiana diferencaEuclidiana_7_6(numero[7][6],20,diff_pixel[7][6]);
	DiferencaEuclidiana diferencaEuclidiana_7_7(numero[7][7],60,diff_pixel[7][7]);
	DiferencaEuclidiana diferencaEuclidiana_7_8(numero[7][8],108,diff_pixel[7][8]);
	DiferencaEuclidiana diferencaEuclidiana_7_9(numero[7][9],125,diff_pixel[7][9]);
	DiferencaEuclidiana diferencaEuclidiana_7_10(numero[7][10],119,diff_pixel[7][10]);
	DiferencaEuclidiana diferencaEuclidiana_8_0(numero[8][0],105,diff_pixel[8][0]);
	DiferencaEuclidiana diferencaEuclidiana_8_1(numero[8][1],131,diff_pixel[8][1]);
	DiferencaEuclidiana diferencaEuclidiana_8_2(numero[8][2],120,diff_pixel[8][2]);
	DiferencaEuclidiana diferencaEuclidiana_8_3(numero[8][3],78,diff_pixel[8][3]);
	DiferencaEuclidiana diferencaEuclidiana_8_4(numero[8][4],28,diff_pixel[8][4]);
	DiferencaEuclidiana diferencaEuclidiana_8_5(numero[8][5],4,diff_pixel[8][5]);
	DiferencaEuclidiana diferencaEuclidiana_8_6(numero[8][6],22,diff_pixel[8][6]);
	DiferencaEuclidiana diferencaEuclidiana_8_7(numero[8][7],62,diff_pixel[8][7]);
	DiferencaEuclidiana diferencaEuclidiana_8_8(numero[8][8],115,diff_pixel[8][8]);
	DiferencaEuclidiana diferencaEuclidiana_8_9(numero[8][9],134,diff_pixel[8][9]);
	DiferencaEuclidiana diferencaEuclidiana_8_10(numero[8][10],118,diff_pixel[8][10]);
	DiferencaEuclidiana diferencaEuclidiana_9_0(numero[9][0],58,diff_pixel[9][0]);
	DiferencaEuclidiana diferencaEuclidiana_9_1(numero[9][1],95,diff_pixel[9][1]);
	DiferencaEuclidiana diferencaEuclidiana_9_2(numero[9][2],131,diff_pixel[9][2]);
	DiferencaEuclidiana diferencaEuclidiana_9_3(numero[9][3],142,diff_pixel[9][3]);
	DiferencaEuclidiana diferencaEuclidiana_9_4(numero[9][4],138,diff_pixel[9][4]);
	DiferencaEuclidiana diferencaEuclidiana_9_5(numero[9][5],134,diff_pixel[9][5]);
	DiferencaEuclidiana diferencaEuclidiana_9_6(numero[9][6],134,diff_pixel[9][6]);
	DiferencaEuclidiana diferencaEuclidiana_9_7(numero[9][7],136,diff_pixel[9][7]);
	DiferencaEuclidiana diferencaEuclidiana_9_8(numero[9][8],134,diff_pixel[9][8]);
	DiferencaEuclidiana diferencaEuclidiana_9_9(numero[9][9],110,diff_pixel[9][9]);
	DiferencaEuclidiana diferencaEuclidiana_9_10(numero[9][10],66,diff_pixel[9][10]);
	DiferencaEuclidiana diferencaEuclidiana_10_0(numero[10][0],16,diff_pixel[10][0]);
	DiferencaEuclidiana diferencaEuclidiana_10_1(numero[10][1],47,diff_pixel[10][1]);
	DiferencaEuclidiana diferencaEuclidiana_10_2(numero[10][2],80,diff_pixel[10][2]);
	DiferencaEuclidiana diferencaEuclidiana_10_3(numero[10][3],103,diff_pixel[10][3]);
	DiferencaEuclidiana diferencaEuclidiana_10_4(numero[10][4],113,diff_pixel[10][4]);
	DiferencaEuclidiana diferencaEuclidiana_10_5(numero[10][5],115,diff_pixel[10][5]);
	DiferencaEuclidiana diferencaEuclidiana_10_6(numero[10][6],119,diff_pixel[10][6]);
	DiferencaEuclidiana diferencaEuclidiana_10_7(numero[10][7],108,diff_pixel[10][7]);
	DiferencaEuclidiana diferencaEuclidiana_10_8(numero[10][8],95,diff_pixel[10][8]);
	DiferencaEuclidiana diferencaEuclidiana_10_9(numero[10][9],64,diff_pixel[10][9]);
	DiferencaEuclidiana diferencaEuclidiana_10_10(numero[10][10],30,diff_pixel[10][10]);
	
endmodule

