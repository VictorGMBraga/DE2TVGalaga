module SomaPixels(
	input [15:0] diff_pixel[3:1][10:0][10:0],
	output [31:0] soma
);

	assign soma =    diff_pixel[1][0][0]
						+ diff_pixel[1][0][1]
						+ diff_pixel[1][0][2]
						+ diff_pixel[1][0][3]
						+ diff_pixel[1][0][4]
						+ diff_pixel[1][0][5]
						+ diff_pixel[1][0][6]
						+ diff_pixel[1][0][7]
						+ diff_pixel[1][0][8]
						+ diff_pixel[1][0][9]
						+ diff_pixel[1][0][10]
						+ diff_pixel[1][1][0]
						+ diff_pixel[1][1][1]
						+ diff_pixel[1][1][2]
						+ diff_pixel[1][1][3]
						+ diff_pixel[1][1][4]
						+ diff_pixel[1][1][5]
						+ diff_pixel[1][1][6]
						+ diff_pixel[1][1][7]
						+ diff_pixel[1][1][8]
						+ diff_pixel[1][1][9]
						+ diff_pixel[1][1][10]
						+ diff_pixel[1][2][0]
						+ diff_pixel[1][2][1]
						+ diff_pixel[1][2][2]
						+ diff_pixel[1][2][3]
						+ diff_pixel[1][2][4]
						+ diff_pixel[1][2][5]
						+ diff_pixel[1][2][6]
						+ diff_pixel[1][2][7]
						+ diff_pixel[1][2][8]
						+ diff_pixel[1][2][9]
						+ diff_pixel[1][2][10]
						+ diff_pixel[1][3][0]
						+ diff_pixel[1][3][1]
						+ diff_pixel[1][3][2]
						+ diff_pixel[1][3][3]
						+ diff_pixel[1][3][4]
						+ diff_pixel[1][3][5]
						+ diff_pixel[1][3][6]
						+ diff_pixel[1][3][7]
						+ diff_pixel[1][3][8]
						+ diff_pixel[1][3][9]
						+ diff_pixel[1][3][10]
						+ diff_pixel[1][4][0]
						+ diff_pixel[1][4][1]
						+ diff_pixel[1][4][2]
						+ diff_pixel[1][4][3]
						+ diff_pixel[1][4][4]
						+ diff_pixel[1][4][5]
						+ diff_pixel[1][4][6]
						+ diff_pixel[1][4][7]
						+ diff_pixel[1][4][8]
						+ diff_pixel[1][4][9]
						+ diff_pixel[1][4][10]
						+ diff_pixel[1][5][0]
						+ diff_pixel[1][5][1]
						+ diff_pixel[1][5][2]
						+ diff_pixel[1][5][3]
						+ diff_pixel[1][5][4]
						+ diff_pixel[1][5][5]
						+ diff_pixel[1][5][6]
						+ diff_pixel[1][5][7]
						+ diff_pixel[1][5][8]
						+ diff_pixel[1][5][9]
						+ diff_pixel[1][5][10]
						+ diff_pixel[1][6][0]
						+ diff_pixel[1][6][1]
						+ diff_pixel[1][6][2]
						+ diff_pixel[1][6][3]
						+ diff_pixel[1][6][4]
						+ diff_pixel[1][6][5]
						+ diff_pixel[1][6][6]
						+ diff_pixel[1][6][7]
						+ diff_pixel[1][6][8]
						+ diff_pixel[1][6][9]
						+ diff_pixel[1][6][10]
						+ diff_pixel[1][7][0]
						+ diff_pixel[1][7][1]
						+ diff_pixel[1][7][2]
						+ diff_pixel[1][7][3]
						+ diff_pixel[1][7][4]
						+ diff_pixel[1][7][5]
						+ diff_pixel[1][7][6]
						+ diff_pixel[1][7][7]
						+ diff_pixel[1][7][8]
						+ diff_pixel[1][7][9]
						+ diff_pixel[1][7][10]
						+ diff_pixel[1][8][0]
						+ diff_pixel[1][8][1]
						+ diff_pixel[1][8][2]
						+ diff_pixel[1][8][3]
						+ diff_pixel[1][8][4]
						+ diff_pixel[1][8][5]
						+ diff_pixel[1][8][6]
						+ diff_pixel[1][8][7]
						+ diff_pixel[1][8][8]
						+ diff_pixel[1][8][9]
						+ diff_pixel[1][8][10]
						+ diff_pixel[1][9][0]
						+ diff_pixel[1][9][1]
						+ diff_pixel[1][9][2]
						+ diff_pixel[1][9][3]
						+ diff_pixel[1][9][4]
						+ diff_pixel[1][9][5]
						+ diff_pixel[1][9][6]
						+ diff_pixel[1][9][7]
						+ diff_pixel[1][9][8]
						+ diff_pixel[1][9][9]
						+ diff_pixel[1][9][10]
						+ diff_pixel[1][10][0]
						+ diff_pixel[1][10][1]
						+ diff_pixel[1][10][2]
						+ diff_pixel[1][10][3]
						+ diff_pixel[1][10][4]
						+ diff_pixel[1][10][5]
						+ diff_pixel[1][10][6]
						+ diff_pixel[1][10][7]
						+ diff_pixel[1][10][8]
						+ diff_pixel[1][10][9]
						+ diff_pixel[1][10][10]
						+ diff_pixel[2][0][0]
						+ diff_pixel[2][0][1]
						+ diff_pixel[2][0][2]
						+ diff_pixel[2][0][3]
						+ diff_pixel[2][0][4]
						+ diff_pixel[2][0][5]
						+ diff_pixel[2][0][6]
						+ diff_pixel[2][0][7]
						+ diff_pixel[2][0][8]
						+ diff_pixel[2][0][9]
						+ diff_pixel[2][0][10]
						+ diff_pixel[2][1][0]
						+ diff_pixel[2][1][1]
						+ diff_pixel[2][1][2]
						+ diff_pixel[2][1][3]
						+ diff_pixel[2][1][4]
						+ diff_pixel[2][1][5]
						+ diff_pixel[2][1][6]
						+ diff_pixel[2][1][7]
						+ diff_pixel[2][1][8]
						+ diff_pixel[2][1][9]
						+ diff_pixel[2][1][10]
						+ diff_pixel[2][2][0]
						+ diff_pixel[2][2][1]
						+ diff_pixel[2][2][2]
						+ diff_pixel[2][2][3]
						+ diff_pixel[2][2][4]
						+ diff_pixel[2][2][5]
						+ diff_pixel[2][2][6]
						+ diff_pixel[2][2][7]
						+ diff_pixel[2][2][8]
						+ diff_pixel[2][2][9]
						+ diff_pixel[2][2][10]
						+ diff_pixel[2][3][0]
						+ diff_pixel[2][3][1]
						+ diff_pixel[2][3][2]
						+ diff_pixel[2][3][3]
						+ diff_pixel[2][3][4]
						+ diff_pixel[2][3][5]
						+ diff_pixel[2][3][6]
						+ diff_pixel[2][3][7]
						+ diff_pixel[2][3][8]
						+ diff_pixel[2][3][9]
						+ diff_pixel[2][3][10]
						+ diff_pixel[2][4][0]
						+ diff_pixel[2][4][1]
						+ diff_pixel[2][4][2]
						+ diff_pixel[2][4][3]
						+ diff_pixel[2][4][4]
						+ diff_pixel[2][4][5]
						+ diff_pixel[2][4][6]
						+ diff_pixel[2][4][7]
						+ diff_pixel[2][4][8]
						+ diff_pixel[2][4][9]
						+ diff_pixel[2][4][10]
						+ diff_pixel[2][5][0]
						+ diff_pixel[2][5][1]
						+ diff_pixel[2][5][2]
						+ diff_pixel[2][5][3]
						+ diff_pixel[2][5][4]
						+ diff_pixel[2][5][5]
						+ diff_pixel[2][5][6]
						+ diff_pixel[2][5][7]
						+ diff_pixel[2][5][8]
						+ diff_pixel[2][5][9]
						+ diff_pixel[2][5][10]
						+ diff_pixel[2][6][0]
						+ diff_pixel[2][6][1]
						+ diff_pixel[2][6][2]
						+ diff_pixel[2][6][3]
						+ diff_pixel[2][6][4]
						+ diff_pixel[2][6][5]
						+ diff_pixel[2][6][6]
						+ diff_pixel[2][6][7]
						+ diff_pixel[2][6][8]
						+ diff_pixel[2][6][9]
						+ diff_pixel[2][6][10]
						+ diff_pixel[2][7][0]
						+ diff_pixel[2][7][1]
						+ diff_pixel[2][7][2]
						+ diff_pixel[2][7][3]
						+ diff_pixel[2][7][4]
						+ diff_pixel[2][7][5]
						+ diff_pixel[2][7][6]
						+ diff_pixel[2][7][7]
						+ diff_pixel[2][7][8]
						+ diff_pixel[2][7][9]
						+ diff_pixel[2][7][10]
						+ diff_pixel[2][8][0]
						+ diff_pixel[2][8][1]
						+ diff_pixel[2][8][2]
						+ diff_pixel[2][8][3]
						+ diff_pixel[2][8][4]
						+ diff_pixel[2][8][5]
						+ diff_pixel[2][8][6]
						+ diff_pixel[2][8][7]
						+ diff_pixel[2][8][8]
						+ diff_pixel[2][8][9]
						+ diff_pixel[2][8][10]
						+ diff_pixel[2][9][0]
						+ diff_pixel[2][9][1]
						+ diff_pixel[2][9][2]
						+ diff_pixel[2][9][3]
						+ diff_pixel[2][9][4]
						+ diff_pixel[2][9][5]
						+ diff_pixel[2][9][6]
						+ diff_pixel[2][9][7]
						+ diff_pixel[2][9][8]
						+ diff_pixel[2][9][9]
						+ diff_pixel[2][9][10]
						+ diff_pixel[2][10][0]
						+ diff_pixel[2][10][1]
						+ diff_pixel[2][10][2]
						+ diff_pixel[2][10][3]
						+ diff_pixel[2][10][4]
						+ diff_pixel[2][10][5]
						+ diff_pixel[2][10][6]
						+ diff_pixel[2][10][7]
						+ diff_pixel[2][10][8]
						+ diff_pixel[2][10][9]
						+ diff_pixel[2][10][10]
						+ diff_pixel[3][0][0]
						+ diff_pixel[3][0][1]
						+ diff_pixel[3][0][2]
						+ diff_pixel[3][0][3]
						+ diff_pixel[3][0][4]
						+ diff_pixel[3][0][5]
						+ diff_pixel[3][0][6]
						+ diff_pixel[3][0][7]
						+ diff_pixel[3][0][8]
						+ diff_pixel[3][0][9]
						+ diff_pixel[3][0][10]
						+ diff_pixel[3][1][0]
						+ diff_pixel[3][1][1]
						+ diff_pixel[3][1][2]
						+ diff_pixel[3][1][3]
						+ diff_pixel[3][1][4]
						+ diff_pixel[3][1][5]
						+ diff_pixel[3][1][6]
						+ diff_pixel[3][1][7]
						+ diff_pixel[3][1][8]
						+ diff_pixel[3][1][9]
						+ diff_pixel[3][1][10]
						+ diff_pixel[3][2][0]
						+ diff_pixel[3][2][1]
						+ diff_pixel[3][2][2]
						+ diff_pixel[3][2][3]
						+ diff_pixel[3][2][4]
						+ diff_pixel[3][2][5]
						+ diff_pixel[3][2][6]
						+ diff_pixel[3][2][7]
						+ diff_pixel[3][2][8]
						+ diff_pixel[3][2][9]
						+ diff_pixel[3][2][10]
						+ diff_pixel[3][3][0]
						+ diff_pixel[3][3][1]
						+ diff_pixel[3][3][2]
						+ diff_pixel[3][3][3]
						+ diff_pixel[3][3][4]
						+ diff_pixel[3][3][5]
						+ diff_pixel[3][3][6]
						+ diff_pixel[3][3][7]
						+ diff_pixel[3][3][8]
						+ diff_pixel[3][3][9]
						+ diff_pixel[3][3][10]
						+ diff_pixel[3][4][0]
						+ diff_pixel[3][4][1]
						+ diff_pixel[3][4][2]
						+ diff_pixel[3][4][3]
						+ diff_pixel[3][4][4]
						+ diff_pixel[3][4][5]
						+ diff_pixel[3][4][6]
						+ diff_pixel[3][4][7]
						+ diff_pixel[3][4][8]
						+ diff_pixel[3][4][9]
						+ diff_pixel[3][4][10]
						+ diff_pixel[3][5][0]
						+ diff_pixel[3][5][1]
						+ diff_pixel[3][5][2]
						+ diff_pixel[3][5][3]
						+ diff_pixel[3][5][4]
						+ diff_pixel[3][5][5]
						+ diff_pixel[3][5][6]
						+ diff_pixel[3][5][7]
						+ diff_pixel[3][5][8]
						+ diff_pixel[3][5][9]
						+ diff_pixel[3][5][10]
						+ diff_pixel[3][6][0]
						+ diff_pixel[3][6][1]
						+ diff_pixel[3][6][2]
						+ diff_pixel[3][6][3]
						+ diff_pixel[3][6][4]
						+ diff_pixel[3][6][5]
						+ diff_pixel[3][6][6]
						+ diff_pixel[3][6][7]
						+ diff_pixel[3][6][8]
						+ diff_pixel[3][6][9]
						+ diff_pixel[3][6][10]
						+ diff_pixel[3][7][0]
						+ diff_pixel[3][7][1]
						+ diff_pixel[3][7][2]
						+ diff_pixel[3][7][3]
						+ diff_pixel[3][7][4]
						+ diff_pixel[3][7][5]
						+ diff_pixel[3][7][6]
						+ diff_pixel[3][7][7]
						+ diff_pixel[3][7][8]
						+ diff_pixel[3][7][9]
						+ diff_pixel[3][7][10]
						+ diff_pixel[3][8][0]
						+ diff_pixel[3][8][1]
						+ diff_pixel[3][8][2]
						+ diff_pixel[3][8][3]
						+ diff_pixel[3][8][4]
						+ diff_pixel[3][8][5]
						+ diff_pixel[3][8][6]
						+ diff_pixel[3][8][7]
						+ diff_pixel[3][8][8]
						+ diff_pixel[3][8][9]
						+ diff_pixel[3][8][10]
						+ diff_pixel[3][9][0]
						+ diff_pixel[3][9][1]
						+ diff_pixel[3][9][2]
						+ diff_pixel[3][9][3]
						+ diff_pixel[3][9][4]
						+ diff_pixel[3][9][5]
						+ diff_pixel[3][9][6]
						+ diff_pixel[3][9][7]
						+ diff_pixel[3][9][8]
						+ diff_pixel[3][9][9]
						+ diff_pixel[3][9][10]
						+ diff_pixel[3][10][0]
						+ diff_pixel[3][10][1]
						+ diff_pixel[3][10][2]
						+ diff_pixel[3][10][3]
						+ diff_pixel[3][10][4]
						+ diff_pixel[3][10][5]
						+ diff_pixel[3][10][6]
						+ diff_pixel[3][10][7]
						+ diff_pixel[3][10][8]
						+ diff_pixel[3][10][9]
						+ diff_pixel[3][10][10];

endmodule
