module SomaPixels(
	input [7:0] diff_pixel[10:0][10:0],
	output [15:0] soma
);

	assign soma =    diff_pixel[0][0]
						+ diff_pixel[0][1]
						+ diff_pixel[0][2]
						+ diff_pixel[0][3]
						+ diff_pixel[0][4]
						+ diff_pixel[0][5]
						+ diff_pixel[0][6]
						+ diff_pixel[0][7]
						+ diff_pixel[0][8]
						+ diff_pixel[0][9]
						+ diff_pixel[0][10]
						+ diff_pixel[1][0]
						+ diff_pixel[1][1]
						+ diff_pixel[1][2]
						+ diff_pixel[1][3]
						+ diff_pixel[1][4]
						+ diff_pixel[1][5]
						+ diff_pixel[1][6]
						+ diff_pixel[1][7]
						+ diff_pixel[1][8]
						+ diff_pixel[1][9]
						+ diff_pixel[1][10]
						+ diff_pixel[2][0]
						+ diff_pixel[2][1]
						+ diff_pixel[2][2]
						+ diff_pixel[2][3]
						+ diff_pixel[2][4]
						+ diff_pixel[2][5]
						+ diff_pixel[2][6]
						+ diff_pixel[2][7]
						+ diff_pixel[2][8]
						+ diff_pixel[2][9]
						+ diff_pixel[2][10]
						+ diff_pixel[3][0]
						+ diff_pixel[3][1]
						+ diff_pixel[3][2]
						+ diff_pixel[3][3]
						+ diff_pixel[3][4]
						+ diff_pixel[3][5]
						+ diff_pixel[3][6]
						+ diff_pixel[3][7]
						+ diff_pixel[3][8]
						+ diff_pixel[3][9]
						+ diff_pixel[3][10]
						+ diff_pixel[4][0]
						+ diff_pixel[4][1]
						+ diff_pixel[4][2]
						+ diff_pixel[4][3]
						+ diff_pixel[4][4]
						+ diff_pixel[4][5]
						+ diff_pixel[4][6]
						+ diff_pixel[4][7]
						+ diff_pixel[4][8]
						+ diff_pixel[4][9]
						+ diff_pixel[4][10]
						+ diff_pixel[5][0]
						+ diff_pixel[5][1]
						+ diff_pixel[5][2]
						+ diff_pixel[5][3]
						+ diff_pixel[5][4]
						+ diff_pixel[5][5]
						+ diff_pixel[5][6]
						+ diff_pixel[5][7]
						+ diff_pixel[5][8]
						+ diff_pixel[5][9]
						+ diff_pixel[5][10]
						+ diff_pixel[6][0]
						+ diff_pixel[6][1]
						+ diff_pixel[6][2]
						+ diff_pixel[6][3]
						+ diff_pixel[6][4]
						+ diff_pixel[6][5]
						+ diff_pixel[6][6]
						+ diff_pixel[6][7]
						+ diff_pixel[6][8]
						+ diff_pixel[6][9]
						+ diff_pixel[6][10]
						+ diff_pixel[7][0]
						+ diff_pixel[7][1]
						+ diff_pixel[7][2]
						+ diff_pixel[7][3]
						+ diff_pixel[7][4]
						+ diff_pixel[7][5]
						+ diff_pixel[7][6]
						+ diff_pixel[7][7]
						+ diff_pixel[7][8]
						+ diff_pixel[7][9]
						+ diff_pixel[7][10]
						+ diff_pixel[8][0]
						+ diff_pixel[8][1]
						+ diff_pixel[8][2]
						+ diff_pixel[8][3]
						+ diff_pixel[8][4]
						+ diff_pixel[8][5]
						+ diff_pixel[8][6]
						+ diff_pixel[8][7]
						+ diff_pixel[8][8]
						+ diff_pixel[8][9]
						+ diff_pixel[8][10]
						+ diff_pixel[9][0]
						+ diff_pixel[9][1]
						+ diff_pixel[9][2]
						+ diff_pixel[9][3]
						+ diff_pixel[9][4]
						+ diff_pixel[9][5]
						+ diff_pixel[9][6]
						+ diff_pixel[9][7]
						+ diff_pixel[9][8]
						+ diff_pixel[9][9]
						+ diff_pixel[9][10]
						+ diff_pixel[10][0]
						+ diff_pixel[10][1]
						+ diff_pixel[10][2]
						+ diff_pixel[10][3]
						+ diff_pixel[10][4]
						+ diff_pixel[10][5]
						+ diff_pixel[10][6]
						+ diff_pixel[10][7]
						+ diff_pixel[10][8]
						+ diff_pixel[10][9]
						+ diff_pixel[10][10];

endmodule
