module Diferenca5(
	input  [7:0] numero[10:0][10:0],
	output [7:0] diff_pixel[10:0][10:0]
);
	
	DiferencaEuclidiana diferencaEuclidiana_00_00(numero[00][00],54,diff_pixel[00][00]);
	DiferencaEuclidiana diferencaEuclidiana_00_01(numero[00][01],80,diff_pixel[00][01]);
	DiferencaEuclidiana diferencaEuclidiana_00_02(numero[00][02],96,diff_pixel[00][02]);
	DiferencaEuclidiana diferencaEuclidiana_00_03(numero[00][03],101,diff_pixel[00][03]);
	DiferencaEuclidiana diferencaEuclidiana_00_04(numero[00][04],98,diff_pixel[00][04]);
	DiferencaEuclidiana diferencaEuclidiana_00_05(numero[00][05],97,diff_pixel[00][05]);
	DiferencaEuclidiana diferencaEuclidiana_00_06(numero[00][06],98,diff_pixel[00][06]);
	DiferencaEuclidiana diferencaEuclidiana_00_07(numero[00][07],91,diff_pixel[00][07]);
	DiferencaEuclidiana diferencaEuclidiana_00_08(numero[00][08],76,diff_pixel[00][08]);
	DiferencaEuclidiana diferencaEuclidiana_00_09(numero[00][09],51,diff_pixel[00][09]);
	DiferencaEuclidiana diferencaEuclidiana_00_10(numero[00][10],22,diff_pixel[00][10]);
	DiferencaEuclidiana diferencaEuclidiana_01_00(numero[01][00],106,diff_pixel[01][00]);
	DiferencaEuclidiana diferencaEuclidiana_01_01(numero[01][01],145,diff_pixel[01][01]);
	DiferencaEuclidiana diferencaEuclidiana_01_02(numero[01][02],164,diff_pixel[01][02]);
	DiferencaEuclidiana diferencaEuclidiana_01_03(numero[01][03],158,diff_pixel[01][03]);
	DiferencaEuclidiana diferencaEuclidiana_01_04(numero[01][04],143,diff_pixel[01][04]);
	DiferencaEuclidiana diferencaEuclidiana_01_05(numero[01][05],135,diff_pixel[01][05]);
	DiferencaEuclidiana diferencaEuclidiana_01_06(numero[01][06],133,diff_pixel[01][06]);
	DiferencaEuclidiana diferencaEuclidiana_01_07(numero[01][07],123,diff_pixel[01][07]);
	DiferencaEuclidiana diferencaEuclidiana_01_08(numero[01][08],104,diff_pixel[01][08]);
	DiferencaEuclidiana diferencaEuclidiana_01_09(numero[01][09],69,diff_pixel[01][09]);
	DiferencaEuclidiana diferencaEuclidiana_01_10(numero[01][10],31,diff_pixel[01][10]);
	DiferencaEuclidiana diferencaEuclidiana_02_00(numero[02][00],106,diff_pixel[02][00]);
	DiferencaEuclidiana diferencaEuclidiana_02_01(numero[02][01],133,diff_pixel[02][01]);
	DiferencaEuclidiana diferencaEuclidiana_02_02(numero[02][02],127,diff_pixel[02][02]);
	DiferencaEuclidiana diferencaEuclidiana_02_03(numero[02][03],86,diff_pixel[02][03]);
	DiferencaEuclidiana diferencaEuclidiana_02_04(numero[02][04],41,diff_pixel[02][04]);
	DiferencaEuclidiana diferencaEuclidiana_02_05(numero[02][05],14,diff_pixel[02][05]);
	DiferencaEuclidiana diferencaEuclidiana_02_06(numero[02][06],2,diff_pixel[02][06]);
	DiferencaEuclidiana diferencaEuclidiana_02_07(numero[02][07],2,diff_pixel[02][07]);
	DiferencaEuclidiana diferencaEuclidiana_02_08(numero[02][08],0,diff_pixel[02][08]);
	DiferencaEuclidiana diferencaEuclidiana_02_09(numero[02][09],0,diff_pixel[02][09]);
	DiferencaEuclidiana diferencaEuclidiana_02_10(numero[02][10],0,diff_pixel[02][10]);
	DiferencaEuclidiana diferencaEuclidiana_03_00(numero[03][00],104,diff_pixel[03][00]);
	DiferencaEuclidiana diferencaEuclidiana_03_01(numero[03][01],143,diff_pixel[03][01]);
	DiferencaEuclidiana diferencaEuclidiana_03_02(numero[03][02],155,diff_pixel[03][02]);
	DiferencaEuclidiana diferencaEuclidiana_03_03(numero[03][03],144,diff_pixel[03][03]);
	DiferencaEuclidiana diferencaEuclidiana_03_04(numero[03][04],125,diff_pixel[03][04]);
	DiferencaEuclidiana diferencaEuclidiana_03_05(numero[03][05],113,diff_pixel[03][05]);
	DiferencaEuclidiana diferencaEuclidiana_03_06(numero[03][06],112,diff_pixel[03][06]);
	DiferencaEuclidiana diferencaEuclidiana_03_07(numero[03][07],105,diff_pixel[03][07]);
	DiferencaEuclidiana diferencaEuclidiana_03_08(numero[03][08],89,diff_pixel[03][08]);
	DiferencaEuclidiana diferencaEuclidiana_03_09(numero[03][09],60,diff_pixel[03][09]);
	DiferencaEuclidiana diferencaEuclidiana_03_10(numero[03][10],33,diff_pixel[03][10]);
	DiferencaEuclidiana diferencaEuclidiana_04_00(numero[04][00],73,diff_pixel[04][00]);
	DiferencaEuclidiana diferencaEuclidiana_04_01(numero[04][01],107,diff_pixel[04][01]);
	DiferencaEuclidiana diferencaEuclidiana_04_02(numero[04][02],122,diff_pixel[04][02]);
	DiferencaEuclidiana diferencaEuclidiana_04_03(numero[04][03],128,diff_pixel[04][03]);
	DiferencaEuclidiana diferencaEuclidiana_04_04(numero[04][04],122,diff_pixel[04][04]);
	DiferencaEuclidiana diferencaEuclidiana_04_05(numero[04][05],123,diff_pixel[04][05]);
	DiferencaEuclidiana diferencaEuclidiana_04_06(numero[04][06],128,diff_pixel[04][06]);
	DiferencaEuclidiana diferencaEuclidiana_04_07(numero[04][07],132,diff_pixel[04][07]);
	DiferencaEuclidiana diferencaEuclidiana_04_08(numero[04][08],123,diff_pixel[04][08]);
	DiferencaEuclidiana diferencaEuclidiana_04_09(numero[04][09],98,diff_pixel[04][09]);
	DiferencaEuclidiana diferencaEuclidiana_04_10(numero[04][10],69,diff_pixel[04][10]);
	DiferencaEuclidiana diferencaEuclidiana_05_00(numero[05][00],0,diff_pixel[05][00]);
	DiferencaEuclidiana diferencaEuclidiana_05_01(numero[05][01],7,diff_pixel[05][01]);
	DiferencaEuclidiana diferencaEuclidiana_05_02(numero[05][02],5,diff_pixel[05][02]);
	DiferencaEuclidiana diferencaEuclidiana_05_03(numero[05][03],6,diff_pixel[05][03]);
	DiferencaEuclidiana diferencaEuclidiana_05_04(numero[05][04],2,diff_pixel[05][04]);
	DiferencaEuclidiana diferencaEuclidiana_05_05(numero[05][05],8,diff_pixel[05][05]);
	DiferencaEuclidiana diferencaEuclidiana_05_06(numero[05][06],29,diff_pixel[05][06]);
	DiferencaEuclidiana diferencaEuclidiana_05_07(numero[05][07],64,diff_pixel[05][07]);
	DiferencaEuclidiana diferencaEuclidiana_05_08(numero[05][08],106,diff_pixel[05][08]);
	DiferencaEuclidiana diferencaEuclidiana_05_09(numero[05][09],118,diff_pixel[05][09]);
	DiferencaEuclidiana diferencaEuclidiana_05_10(numero[05][10],120,diff_pixel[05][10]);
	DiferencaEuclidiana diferencaEuclidiana_06_00(numero[06][00],1,diff_pixel[06][00]);
	DiferencaEuclidiana diferencaEuclidiana_06_01(numero[06][01],0,diff_pixel[06][01]);
	DiferencaEuclidiana diferencaEuclidiana_06_02(numero[06][02],0,diff_pixel[06][02]);
	DiferencaEuclidiana diferencaEuclidiana_06_03(numero[06][03],0,diff_pixel[06][03]);
	DiferencaEuclidiana diferencaEuclidiana_06_04(numero[06][04],0,diff_pixel[06][04]);
	DiferencaEuclidiana diferencaEuclidiana_06_05(numero[06][05],0,diff_pixel[06][05]);
	DiferencaEuclidiana diferencaEuclidiana_06_06(numero[06][06],24,diff_pixel[06][06]);
	DiferencaEuclidiana diferencaEuclidiana_06_07(numero[06][07],61,diff_pixel[06][07]);
	DiferencaEuclidiana diferencaEuclidiana_06_08(numero[06][08],109,diff_pixel[06][08]);
	DiferencaEuclidiana diferencaEuclidiana_06_09(numero[06][09],126,diff_pixel[06][09]);
	DiferencaEuclidiana diferencaEuclidiana_06_10(numero[06][10],125,diff_pixel[06][10]);
	DiferencaEuclidiana diferencaEuclidiana_07_00(numero[07][00],42,diff_pixel[07][00]);
	DiferencaEuclidiana diferencaEuclidiana_07_01(numero[07][01],37,diff_pixel[07][01]);
	DiferencaEuclidiana diferencaEuclidiana_07_02(numero[07][02],31,diff_pixel[07][02]);
	DiferencaEuclidiana diferencaEuclidiana_07_03(numero[07][03],19,diff_pixel[07][03]);
	DiferencaEuclidiana diferencaEuclidiana_07_04(numero[07][04],3,diff_pixel[07][04]);
	DiferencaEuclidiana diferencaEuclidiana_07_05(numero[07][05],0,diff_pixel[07][05]);
	DiferencaEuclidiana diferencaEuclidiana_07_06(numero[07][06],22,diff_pixel[07][06]);
	DiferencaEuclidiana diferencaEuclidiana_07_07(numero[07][07],59,diff_pixel[07][07]);
	DiferencaEuclidiana diferencaEuclidiana_07_08(numero[07][08],106,diff_pixel[07][08]);
	DiferencaEuclidiana diferencaEuclidiana_07_09(numero[07][09],122,diff_pixel[07][09]);
	DiferencaEuclidiana diferencaEuclidiana_07_10(numero[07][10],120,diff_pixel[07][10]);
	DiferencaEuclidiana diferencaEuclidiana_08_00(numero[08][00],99,diff_pixel[08][00]);
	DiferencaEuclidiana diferencaEuclidiana_08_01(numero[08][01],125,diff_pixel[08][01]);
	DiferencaEuclidiana diferencaEuclidiana_08_02(numero[08][02],120,diff_pixel[08][02]);
	DiferencaEuclidiana diferencaEuclidiana_08_03(numero[08][03],78,diff_pixel[08][03]);
	DiferencaEuclidiana diferencaEuclidiana_08_04(numero[08][04],28,diff_pixel[08][04]);
	DiferencaEuclidiana diferencaEuclidiana_08_05(numero[08][05],4,diff_pixel[08][05]);
	DiferencaEuclidiana diferencaEuclidiana_08_06(numero[08][06],21,diff_pixel[08][06]);
	DiferencaEuclidiana diferencaEuclidiana_08_07(numero[08][07],61,diff_pixel[08][07]);
	DiferencaEuclidiana diferencaEuclidiana_08_08(numero[08][08],116,diff_pixel[08][08]);
	DiferencaEuclidiana diferencaEuclidiana_08_09(numero[08][09],133,diff_pixel[08][09]);
	DiferencaEuclidiana diferencaEuclidiana_08_10(numero[08][10],121,diff_pixel[08][10]);
	DiferencaEuclidiana diferencaEuclidiana_09_00(numero[09][00],52,diff_pixel[09][00]);
	DiferencaEuclidiana diferencaEuclidiana_09_01(numero[09][01],92,diff_pixel[09][01]);
	DiferencaEuclidiana diferencaEuclidiana_09_02(numero[09][02],131,diff_pixel[09][02]);
	DiferencaEuclidiana diferencaEuclidiana_09_03(numero[09][03],139,diff_pixel[09][03]);
	DiferencaEuclidiana diferencaEuclidiana_09_04(numero[09][04],137,diff_pixel[09][04]);
	DiferencaEuclidiana diferencaEuclidiana_09_05(numero[09][05],132,diff_pixel[09][05]);
	DiferencaEuclidiana diferencaEuclidiana_09_06(numero[09][06],134,diff_pixel[09][06]);
	DiferencaEuclidiana diferencaEuclidiana_09_07(numero[09][07],136,diff_pixel[09][07]);
	DiferencaEuclidiana diferencaEuclidiana_09_08(numero[09][08],134,diff_pixel[09][08]);
	DiferencaEuclidiana diferencaEuclidiana_09_09(numero[09][09],109,diff_pixel[09][09]);
	DiferencaEuclidiana diferencaEuclidiana_09_10(numero[09][10],67,diff_pixel[09][10]);
	DiferencaEuclidiana diferencaEuclidiana_10_00(numero[10][00],15,diff_pixel[10][00]);
	DiferencaEuclidiana diferencaEuclidiana_10_01(numero[10][01],47,diff_pixel[10][01]);
	DiferencaEuclidiana diferencaEuclidiana_10_02(numero[10][02],82,diff_pixel[10][02]);
	DiferencaEuclidiana diferencaEuclidiana_10_03(numero[10][03],105,diff_pixel[10][03]);
	DiferencaEuclidiana diferencaEuclidiana_10_04(numero[10][04],115,diff_pixel[10][04]);
	DiferencaEuclidiana diferencaEuclidiana_10_05(numero[10][05],116,diff_pixel[10][05]);
	DiferencaEuclidiana diferencaEuclidiana_10_06(numero[10][06],119,diff_pixel[10][06]);
	DiferencaEuclidiana diferencaEuclidiana_10_07(numero[10][07],108,diff_pixel[10][07]);
	DiferencaEuclidiana diferencaEuclidiana_10_08(numero[10][08],95,diff_pixel[10][08]);
	DiferencaEuclidiana diferencaEuclidiana_10_09(numero[10][09],64,diff_pixel[10][09]);
	DiferencaEuclidiana diferencaEuclidiana_10_10(numero[10][10],30,diff_pixel[10][10]);	

endmodule
