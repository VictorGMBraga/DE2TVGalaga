module Diferenca2(
	input  [7:0] numero[10:0][10:0],
	output [7:0] diff_pixel[10:0][10:0]
);
	
	DiferencaEuclidiana diferencaEuclidiana_00_00(numero[00][00],30,diff_pixel[00][00]);
	DiferencaEuclidiana diferencaEuclidiana_00_01(numero[00][01],58,diff_pixel[00][01]);
	DiferencaEuclidiana diferencaEuclidiana_00_02(numero[00][02],80,diff_pixel[00][02]);
	DiferencaEuclidiana diferencaEuclidiana_00_03(numero[00][03],101,diff_pixel[00][03]);
	DiferencaEuclidiana diferencaEuclidiana_00_04(numero[00][04],101,diff_pixel[00][04]);
	DiferencaEuclidiana diferencaEuclidiana_00_05(numero[00][05],103,diff_pixel[00][05]);
	DiferencaEuclidiana diferencaEuclidiana_00_06(numero[00][06],99,diff_pixel[00][06]);
	DiferencaEuclidiana diferencaEuclidiana_00_07(numero[00][07],92,diff_pixel[00][07]);
	DiferencaEuclidiana diferencaEuclidiana_00_08(numero[00][08],76,diff_pixel[00][08]);
	DiferencaEuclidiana diferencaEuclidiana_00_09(numero[00][09],51,diff_pixel[00][09]);
	DiferencaEuclidiana diferencaEuclidiana_00_10(numero[00][10],22,diff_pixel[00][10]);
	DiferencaEuclidiana diferencaEuclidiana_01_00(numero[01][00],46,diff_pixel[01][00]);
	DiferencaEuclidiana diferencaEuclidiana_01_01(numero[01][01],89,diff_pixel[01][01]);
	DiferencaEuclidiana diferencaEuclidiana_01_02(numero[01][02],126,diff_pixel[01][02]);
	DiferencaEuclidiana diferencaEuclidiana_01_03(numero[01][03],143,diff_pixel[01][03]);
	DiferencaEuclidiana diferencaEuclidiana_01_04(numero[01][04],143,diff_pixel[01][04]);
	DiferencaEuclidiana diferencaEuclidiana_01_05(numero[01][05],138,diff_pixel[01][05]);
	DiferencaEuclidiana diferencaEuclidiana_01_06(numero[01][06],142,diff_pixel[01][06]);
	DiferencaEuclidiana diferencaEuclidiana_01_07(numero[01][07],140,diff_pixel[01][07]);
	DiferencaEuclidiana diferencaEuclidiana_01_08(numero[01][08],135,diff_pixel[01][08]);
	DiferencaEuclidiana diferencaEuclidiana_01_09(numero[01][09],107,diff_pixel[01][09]);
	DiferencaEuclidiana diferencaEuclidiana_01_10(numero[01][10],62,diff_pixel[01][10]);
	DiferencaEuclidiana diferencaEuclidiana_02_00(numero[02][00],98,diff_pixel[02][00]);
	DiferencaEuclidiana diferencaEuclidiana_02_01(numero[02][01],123,diff_pixel[02][01]);
	DiferencaEuclidiana diferencaEuclidiana_02_02(numero[02][02],117,diff_pixel[02][02]);
	DiferencaEuclidiana diferencaEuclidiana_02_03(numero[02][03],80,diff_pixel[02][03]);
	DiferencaEuclidiana diferencaEuclidiana_02_04(numero[02][04],31,diff_pixel[02][04]);
	DiferencaEuclidiana diferencaEuclidiana_02_05(numero[02][05],9,diff_pixel[02][05]);
	DiferencaEuclidiana diferencaEuclidiana_02_06(numero[02][06],23,diff_pixel[02][06]);
	DiferencaEuclidiana diferencaEuclidiana_02_07(numero[02][07],60,diff_pixel[02][07]);
	DiferencaEuclidiana diferencaEuclidiana_02_08(numero[02][08],107,diff_pixel[02][08]);
	DiferencaEuclidiana diferencaEuclidiana_02_09(numero[02][09],125,diff_pixel[02][09]);
	DiferencaEuclidiana diferencaEuclidiana_02_10(numero[02][10],114,diff_pixel[02][10]);
	DiferencaEuclidiana diferencaEuclidiana_03_00(numero[03][00],31,diff_pixel[03][00]);
	DiferencaEuclidiana diferencaEuclidiana_03_01(numero[03][01],43,diff_pixel[03][01]);
	DiferencaEuclidiana diferencaEuclidiana_03_02(numero[03][02],38,diff_pixel[03][02]);
	DiferencaEuclidiana diferencaEuclidiana_03_03(numero[03][03],21,diff_pixel[03][03]);
	DiferencaEuclidiana diferencaEuclidiana_03_04(numero[03][04],9,diff_pixel[03][04]);
	DiferencaEuclidiana diferencaEuclidiana_03_05(numero[03][05],18,diff_pixel[03][05]);
	DiferencaEuclidiana diferencaEuclidiana_03_06(numero[03][06],54,diff_pixel[03][06]);
	DiferencaEuclidiana diferencaEuclidiana_03_07(numero[03][07],101,diff_pixel[03][07]);
	DiferencaEuclidiana diferencaEuclidiana_03_08(numero[03][08],141,diff_pixel[03][08]);
	DiferencaEuclidiana diferencaEuclidiana_03_09(numero[03][09],142,diff_pixel[03][09]);
	DiferencaEuclidiana diferencaEuclidiana_03_10(numero[03][10],126,diff_pixel[03][10]);
	DiferencaEuclidiana diferencaEuclidiana_04_00(numero[04][00],0,diff_pixel[04][00]);
	DiferencaEuclidiana diferencaEuclidiana_04_01(numero[04][01],0,diff_pixel[04][01]);
	DiferencaEuclidiana diferencaEuclidiana_04_02(numero[04][02],6,diff_pixel[04][02]);
	DiferencaEuclidiana diferencaEuclidiana_04_03(numero[04][03],22,diff_pixel[04][03]);
	DiferencaEuclidiana diferencaEuclidiana_04_04(numero[04][04],48,diff_pixel[04][04]);
	DiferencaEuclidiana diferencaEuclidiana_04_05(numero[04][05],76,diff_pixel[04][05]);
	DiferencaEuclidiana diferencaEuclidiana_04_06(numero[04][06],116,diff_pixel[04][06]);
	DiferencaEuclidiana diferencaEuclidiana_04_07(numero[04][07],146,diff_pixel[04][07]);
	DiferencaEuclidiana diferencaEuclidiana_04_08(numero[04][08],160,diff_pixel[04][08]);
	DiferencaEuclidiana diferencaEuclidiana_04_09(numero[04][09],139,diff_pixel[04][09]);
	DiferencaEuclidiana diferencaEuclidiana_04_10(numero[04][10],114,diff_pixel[04][10]);
	DiferencaEuclidiana diferencaEuclidiana_05_00(numero[05][00],8,diff_pixel[05][00]);
	DiferencaEuclidiana diferencaEuclidiana_05_01(numero[05][01],10,diff_pixel[05][01]);
	DiferencaEuclidiana diferencaEuclidiana_05_02(numero[05][02],39,diff_pixel[05][02]);
	DiferencaEuclidiana diferencaEuclidiana_05_03(numero[05][03],89,diff_pixel[05][03]);
	DiferencaEuclidiana diferencaEuclidiana_05_04(numero[05][04],133,diff_pixel[05][04]);
	DiferencaEuclidiana diferencaEuclidiana_05_05(numero[05][05],159,diff_pixel[05][05]);
	DiferencaEuclidiana diferencaEuclidiana_05_06(numero[05][06],179,diff_pixel[05][06]);
	DiferencaEuclidiana diferencaEuclidiana_05_07(numero[05][07],169,diff_pixel[05][07]);
	DiferencaEuclidiana diferencaEuclidiana_05_08(numero[05][08],145,diff_pixel[05][08]);
	DiferencaEuclidiana diferencaEuclidiana_05_09(numero[05][09],102,diff_pixel[05][09]);
	DiferencaEuclidiana diferencaEuclidiana_05_10(numero[05][10],63,diff_pixel[05][10]);
	DiferencaEuclidiana diferencaEuclidiana_06_00(numero[06][00],26,diff_pixel[06][00]);
	DiferencaEuclidiana diferencaEuclidiana_06_01(numero[06][01],44,diff_pixel[06][01]);
	DiferencaEuclidiana diferencaEuclidiana_06_02(numero[06][02],92,diff_pixel[06][02]);
	DiferencaEuclidiana diferencaEuclidiana_06_03(numero[06][03],138,diff_pixel[06][03]);
	DiferencaEuclidiana diferencaEuclidiana_06_04(numero[06][04],170,diff_pixel[06][04]);
	DiferencaEuclidiana diferencaEuclidiana_06_05(numero[06][05],177,diff_pixel[06][05]);
	DiferencaEuclidiana diferencaEuclidiana_06_06(numero[06][06],167,diff_pixel[06][06]);
	DiferencaEuclidiana diferencaEuclidiana_06_07(numero[06][07],138,diff_pixel[06][07]);
	DiferencaEuclidiana diferencaEuclidiana_06_08(numero[06][08],93,diff_pixel[06][08]);
	DiferencaEuclidiana diferencaEuclidiana_06_09(numero[06][09],50,diff_pixel[06][09]);
	DiferencaEuclidiana diferencaEuclidiana_06_10(numero[06][10],24,diff_pixel[06][10]);
	DiferencaEuclidiana diferencaEuclidiana_07_00(numero[07][00],62,diff_pixel[07][00]);
	DiferencaEuclidiana diferencaEuclidiana_07_01(numero[07][01],89,diff_pixel[07][01]);
	DiferencaEuclidiana diferencaEuclidiana_07_02(numero[07][02],132,diff_pixel[07][02]);
	DiferencaEuclidiana diferencaEuclidiana_07_03(numero[07][03],156,diff_pixel[07][03]);
	DiferencaEuclidiana diferencaEuclidiana_07_04(numero[07][04],159,diff_pixel[07][04]);
	DiferencaEuclidiana diferencaEuclidiana_07_05(numero[07][05],139,diff_pixel[07][05]);
	DiferencaEuclidiana diferencaEuclidiana_07_06(numero[07][06],111,diff_pixel[07][06]);
	DiferencaEuclidiana diferencaEuclidiana_07_07(numero[07][07],79,diff_pixel[07][07]);
	DiferencaEuclidiana diferencaEuclidiana_07_08(numero[07][08],44,diff_pixel[07][08]);
	DiferencaEuclidiana diferencaEuclidiana_07_09(numero[07][09],15,diff_pixel[07][09]);
	DiferencaEuclidiana diferencaEuclidiana_07_10(numero[07][10],5,diff_pixel[07][10]);
	DiferencaEuclidiana diferencaEuclidiana_08_00(numero[08][00],123,diff_pixel[08][00]);
	DiferencaEuclidiana diferencaEuclidiana_08_01(numero[08][01],151,diff_pixel[08][01]);
	DiferencaEuclidiana diferencaEuclidiana_08_02(numero[08][02],166,diff_pixel[08][02]);
	DiferencaEuclidiana diferencaEuclidiana_08_03(numero[08][03],153,diff_pixel[08][03]);
	DiferencaEuclidiana diferencaEuclidiana_08_04(numero[08][04],109,diff_pixel[08][04]);
	DiferencaEuclidiana diferencaEuclidiana_08_05(numero[08][05],52,diff_pixel[08][05]);
	DiferencaEuclidiana diferencaEuclidiana_08_06(numero[08][06],11,diff_pixel[08][06]);
	DiferencaEuclidiana diferencaEuclidiana_08_07(numero[08][07],0,diff_pixel[08][07]);
	DiferencaEuclidiana diferencaEuclidiana_08_08(numero[08][08],0,diff_pixel[08][08]);
	DiferencaEuclidiana diferencaEuclidiana_08_09(numero[08][09],0,diff_pixel[08][09]);
	DiferencaEuclidiana diferencaEuclidiana_08_10(numero[08][10],0,diff_pixel[08][10]);
	DiferencaEuclidiana diferencaEuclidiana_09_00(numero[09][00],106,diff_pixel[09][00]);
	DiferencaEuclidiana diferencaEuclidiana_09_01(numero[09][01],149,diff_pixel[09][01]);
	DiferencaEuclidiana diferencaEuclidiana_09_02(numero[09][02],173,diff_pixel[09][02]);
	DiferencaEuclidiana diferencaEuclidiana_09_03(numero[09][03],175,diff_pixel[09][03]);
	DiferencaEuclidiana diferencaEuclidiana_09_04(numero[09][04],161,diff_pixel[09][04]);
	DiferencaEuclidiana diferencaEuclidiana_09_05(numero[09][05],142,diff_pixel[09][05]);
	DiferencaEuclidiana diferencaEuclidiana_09_06(numero[09][06],129,diff_pixel[09][06]);
	DiferencaEuclidiana diferencaEuclidiana_09_07(numero[09][07],123,diff_pixel[09][07]);
	DiferencaEuclidiana diferencaEuclidiana_09_08(numero[09][08],118,diff_pixel[09][08]);
	DiferencaEuclidiana diferencaEuclidiana_09_09(numero[09][09],104,diff_pixel[09][09]);
	DiferencaEuclidiana diferencaEuclidiana_09_10(numero[09][10],79,diff_pixel[09][10]);
	DiferencaEuclidiana diferencaEuclidiana_10_00(numero[10][00],68,diff_pixel[10][00]);
	DiferencaEuclidiana diferencaEuclidiana_10_01(numero[10][01],103,diff_pixel[10][01]);
	DiferencaEuclidiana diferencaEuclidiana_10_02(numero[10][02],118,diff_pixel[10][02]);
	DiferencaEuclidiana diferencaEuclidiana_10_03(numero[10][03],125,diff_pixel[10][03]);
	DiferencaEuclidiana diferencaEuclidiana_10_04(numero[10][04],121,diff_pixel[10][04]);
	DiferencaEuclidiana diferencaEuclidiana_10_05(numero[10][05],120,diff_pixel[10][05]);
	DiferencaEuclidiana diferencaEuclidiana_10_06(numero[10][06],120,diff_pixel[10][06]);
	DiferencaEuclidiana diferencaEuclidiana_10_07(numero[10][07],121,diff_pixel[10][07]);
	DiferencaEuclidiana diferencaEuclidiana_10_08(numero[10][08],116,diff_pixel[10][08]);
	DiferencaEuclidiana diferencaEuclidiana_10_09(numero[10][09],100,diff_pixel[10][09]);
	DiferencaEuclidiana diferencaEuclidiana_10_10(numero[10][10],80,diff_pixel[10][10]);
	
endmodule

